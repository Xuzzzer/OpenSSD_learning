
`define		D_CPLD_FMT					3'b010
`define		D_CPLD_TYPE					5'b01010
`define		D_CPLD_TC					3'b000
`define		D_CPLD_ATTR1				1'b0
`define		D_CPLD_TH					1'b0
`define		D_CPLD_TD					1'b0
`define		D_CPLD_EP					1'b0
`define		D_CPLD_ATTR2				2'b00
`define		D_CPLD_AT					2'b00
`define		D_CPLD_CS					3'b000
`define		D_CPLD_BCM					1'b0

`define		D_MRD_FMT					3'b001
`define		D_MRD_TYPE					5'b00000
`define		D_MRD_TC					3'b000
`define		D_MRD_ATTR1					1'b0
`define		D_MRD_TH					1'b0
`define		D_MRD_TD					1'b0
`define		D_MRD_EP					1'b0
`define		D_MRD_ATTR2					2'b00
`define		D_MRD_AT					2'b00
`define		D_MRD_LAST_BE				8'b00001111
`define		D_MRD_1ST_BE				8'b00001111

`define		D_MWR_FMT					3'b011
`define		D_MWR_TYPE					5'b00000
`define		D_MWR_TC					3'b000
`define		D_MWR_ATTR1					1'b0
`define		D_MWR_TH					1'b0
`define		D_MWR_TD					1'b0
`define		D_MWR_EP					1'b0
`define		D_MWR_ATTR2					2'b00
`define		D_MWR_AT					2'b00
`define		D_MWR_LAST_BE				8'b00001111
`define		D_MWR_1ST_BE				8'b00001111
