

//   - minor modification for releasing
//
// * v1.1.1
//   - bug fix: state machine
//
// * v1.1.0
//   - change state machine: divide states
//   - insert additional registers
//   - improve frequency characteristic
//
// * v1.0.0
//   - first draft
//   - KES: binary version of inversion-less Berlekamp-Massey algorithm (iBM.b)
//////////////////////////////////////////////////////////////////////////////////

`include "d_KES_parameters.vh"
`timescale 1ns / 1ps

module d_BCH_KES_top
(
	input  wire 						i_clk,
	input  wire 						i_RESET,
	input  wire							i_stop_dec,
    
    input  wire [3:0]                   i_channel_sel,
	input  wire 						i_execute_kes,
    input  wire                         i_data_fowarding,
	input  wire							i_buf_available,
					
	input  wire	     					i_chunk_number,
	input  wire							i_buf_sequence_end,
					
	output reg							o_kes_sequence_end,
	output wire							o_kes_fail,
	output wire							o_kes_available,
	output reg  [3:0]                   o_channel_sel,				
	output reg 	     					o_chunk_number,
	output reg							o_buf_sequence_end,
	
	output reg	[`D_KES_ECC_T_BIT-1:0]	o_error_count,
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// input port: syndrome
	// output port: error locator polynomial term
	
	// syndrome: 63, 2t-1
	// elpt: 33, t+1
	
    input wire [`D_KES_GF_ORDER*(`D_KES_ECC_T*2-1)-1:0] i_syndromes,

    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_000,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_001,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_002,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_003,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_004,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_005,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_006,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_007,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_008,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_009,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_010,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_011,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_012,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_013,
    output wire [`D_KES_GF_ORDER-1:0] 	o_v_2i_014
	
	                                          ///
	                                        /////	
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
);
	
	parameter [11:0] D_KES_VALUE_ZERO = 12'b0000_0000_0000;
	parameter [11:0] D_KES_VALUE_ONE = 12'b0000_0000_0001;
	
	// FSM parameters
	parameter KES_FSM_BIT = 7;
	parameter KES_RESET = 7'b0000001; // reset: w_RESET_KES <= 0
	parameter KES_START = 7'b0000010; // start: SDR capture, w_RESET_KES <= 1
	parameter KES_STEP1 = 7'b0000100; 
	parameter KES_STEP2 = 7'b0001000; 
    parameter KES_FWD   = 7'b0010000;
    parameter KES_PAUSE = 7'b0100000;
	parameter KES_OUT	= 7'b1000000;
	
	
	// variable declaration
	
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// internal wires for PE
	// coef: (1+S)V, v_2i, deg 0 chk bit
	
	// coef: (1+S)V: 33, t+1
	// v_2i: 33, t+1
	// deg 0 chk bit: 34, t+2
	
	wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_000;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_001;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_002;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_003;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_004;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_005;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_006;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_007;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_008;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_009;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_010;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_011;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_012;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_013;
    wire [`D_KES_GF_ORDER-1:0] w_coef_2ip1_014;

    wire w_v_2i_X_deg_chk_bit_000; // from PE_ELU_MINodr
    wire w_v_2i_X_deg_chk_bit_001; // from PE_ELU_sMINodr
    wire w_v_2i_X_deg_chk_bit_002; // from PE_ELU_NMLodr
    wire w_v_2i_X_deg_chk_bit_003; // from PE_ELU_NMLodr
    wire w_v_2i_X_deg_chk_bit_004; // from PE_ELU_NMLodr
    wire w_v_2i_X_deg_chk_bit_005; // from PE_ELU_NMLodr
    wire w_v_2i_X_deg_chk_bit_006; // from PE_ELU_NMLodr
    wire w_v_2i_X_deg_chk_bit_007; // from PE_ELU_NMLodr
    wire w_v_2i_X_deg_chk_bit_008; // from PE_ELU_NMLodr
    wire w_v_2i_X_deg_chk_bit_009; // from PE_ELU_NMLodr
    wire w_v_2i_X_deg_chk_bit_010; // from PE_ELU_NMLodr
    wire w_v_2i_X_deg_chk_bit_011; // from PE_ELU_NMLodr
    wire w_v_2i_X_deg_chk_bit_012; // from PE_ELU_NMLodr
    wire w_v_2i_X_deg_chk_bit_013; // from PE_ELU_NMLodr
    wire w_v_2i_X_deg_chk_bit_014; // from PE_ELU_NMLodr
    wire w_v_2i_X_deg_chk_bit_015; // from PE_ELU_NMLodr
	
	                                          ///
	                                        /////	
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
	
	// registered input
	reg [(`D_KES_ECC_T*2*`D_KES_GF_ORDER)-1:0] r_sdr_buffer;
	
	// encoder FSM state
	reg [KES_FSM_BIT-1:0] r_cur_state;
	reg [KES_FSM_BIT-1:0] r_nxt_state;
	
	reg [`D_KES_L_CNT_BIT-1:0] r_count_kes; // internal counter
	
	reg  r_RESET_kes_sequence;
	wire w_RESET_KES;
	
	wire w_last_interation;
	wire [`D_KES_ECC_T:0]	w_v_error;
	
	wire                       w_d_2i_ZERO_chk_bit;
    wire [`D_KES_GF_ORDER-1:0] w_d_2i;
	
	wire [`D_KES_GF_ORDER-1:0] w_delta_2i;
	reg  [`D_KES_GF_ORDER-1:0] r_delta_2im2;
	reg  [`D_KES_GF_ORDER-1:0] r_delta_2im2_d0; // duplicate register
	
	wire w_condition_2i;
	
	reg r_EXECUTE_PE_DC;
	
	reg r_EXECUTE_PE_ELU;
	
	wire [`D_KES_ECC_T+1:0] w_v_2ip2_deg_info;
	reg  [`D_KES_ECC_T+1:0] r_v_2i_X_deg_chk_bit_b;
	
	
	reg r_ELP_degree_condition_violation;
	reg [`D_KES_ECC_T_BIT-1:0] r_v_2i_maximum_deg;
	reg r_v_2i_deg_condition;
	
	wire [`D_KES_GF_ORDER-1:0] w_sdr_to_DC_001;
	wire [`D_KES_GF_ORDER-1:0] w_sdr_to_DC_000;
	
	reg						   r_buf_sequence_end;
    reg                        r_data_fowarding;
	
	// generate control/indicate signal
	
	assign w_RESET_KES = (i_RESET) | (r_RESET_kes_sequence);	
	
	assign w_last_interation = (r_count_kes == `D_KES_L_CNT);
	assign o_kes_fail = (o_error_count == 4'b1110);
	assign o_kes_available = (r_cur_state == KES_RESET); //|| ((r_cur_state == KES_STEP7) && (o_kes_sequence_end));
	
	assign w_delta_2i[`D_KES_GF_ORDER-1:0] = (w_condition_2i)? (w_d_2i[`D_KES_GF_ORDER-1:0]):(r_delta_2im2[`D_KES_GF_ORDER-1:0]);
	assign w_v_error[`D_KES_ECC_T:0] = { (|o_v_2i_000[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_001[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_002[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_003[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_004[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_005[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_006[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_007[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_008[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_009[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_010[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_011[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_012[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_013[`D_KES_GF_ORDER-1:0]) , (|o_v_2i_014[`D_KES_GF_ORDER-1:0]) };

    assign w_d_2i = w_coef_2ip1_000[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_001[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_002[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_003[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_004[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_005[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_006[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_007[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_008[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_009[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_010[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_011[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_012[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_013[`D_KES_GF_ORDER-1:0]^ w_coef_2ip1_014[`D_KES_GF_ORDER-1:0] ;
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// w_v_2ip2_deg_info
		
	// all deg info: 34, t+2
	
    assign w_v_2ip2_deg_info[`D_KES_ECC_T+1:0] = { w_v_2i_X_deg_chk_bit_015, w_v_2i_X_deg_chk_bit_014, w_v_2i_X_deg_chk_bit_013, w_v_2i_X_deg_chk_bit_012, w_v_2i_X_deg_chk_bit_011, w_v_2i_X_deg_chk_bit_010, w_v_2i_X_deg_chk_bit_009, w_v_2i_X_deg_chk_bit_008, w_v_2i_X_deg_chk_bit_007, w_v_2i_X_deg_chk_bit_006, w_v_2i_X_deg_chk_bit_005, w_v_2i_X_deg_chk_bit_004, w_v_2i_X_deg_chk_bit_003, w_v_2i_X_deg_chk_bit_002, w_v_2i_X_deg_chk_bit_001, w_v_2i_X_deg_chk_bit_000};
	
	                                          ///
	                                        /////	
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
	
	assign w_d_2i_ZERO_chk_bit = |(w_d_2i[`D_KES_GF_ORDER-1:0]);
	always @ ( r_v_2i_maximum_deg, r_count_kes )
	begin	
		// if you change something, handle follow codes carefully
		if ( r_v_2i_maximum_deg > r_count_kes )	begin
			r_v_2i_deg_condition <= 1'b0;
		end	else begin
			r_v_2i_deg_condition <= 1'b1;
		end
	end
	assign w_condition_2i = (w_d_2i_ZERO_chk_bit) & (r_v_2i_deg_condition);
		
	assign w_sdr_to_DC_001[`D_KES_GF_ORDER-1:0] = r_sdr_buffer[(`D_KES_ECC_T*2  )*`D_KES_GF_ORDER-1:(`D_KES_ECC_T*2-1)*`D_KES_GF_ORDER];
	assign w_sdr_to_DC_000[`D_KES_GF_ORDER-1:0] = r_sdr_buffer[(`D_KES_ECC_T*2-1)*`D_KES_GF_ORDER-1:(`D_KES_ECC_T*2-2)*`D_KES_GF_ORDER];
	
	
	
	//FSM
	// update current state to next state
	always @ (posedge i_clk)
	begin
		if ((i_RESET) || (i_stop_dec)) begin
			r_cur_state <= KES_RESET;
		end else begin
			r_cur_state <= r_nxt_state;
		end
	end
	
	// decide next state
	always @ ( * )
	begin
		if (o_kes_fail) begin
			r_nxt_state <= KES_RESET;
		end	else begin
			case (r_cur_state)
			KES_RESET: begin
				r_nxt_state <= (i_execute_kes)? KES_START:KES_RESET;
			end
			KES_START: begin
				r_nxt_state <= (r_data_fowarding)? KES_FWD:KES_STEP1;
			end
			KES_STEP1: begin
				r_nxt_state <= KES_STEP2;
			end
			KES_STEP2: begin
				r_nxt_state <= (w_last_interation)? ((i_buf_available)? (KES_OUT): (KES_PAUSE)):(KES_STEP1);
			end
            KES_FWD: begin
                r_nxt_state <= (i_buf_available)? (KES_OUT): (KES_FWD);
            end
            KES_PAUSE: begin
                r_nxt_state <= (i_buf_available)? (KES_OUT): (KES_PAUSE);
            end
			KES_OUT: begin
				r_nxt_state <= KES_RESET;
			end
			default: begin
				r_nxt_state <= KES_RESET;
			end
			endcase
		end
	end

	// state behaviour
	always @ (posedge i_clk)
	begin
		if ((i_RESET) || (i_stop_dec)) 
			o_kes_sequence_end <= 0;
		else begin
			case (r_nxt_state)
			KES_OUT: 
				o_kes_sequence_end <= 1'b1;
			default: 
				o_kes_sequence_end <= 0;
			endcase
			end
	end
	
	always @ (posedge i_clk)
	begin
		if ((i_RESET) || (i_stop_dec)) begin
			r_count_kes <= 0;
			r_sdr_buffer[(`D_KES_ECC_T*2*`D_KES_GF_ORDER)-1:0] <= 0;
			r_RESET_kes_sequence <= 1;
			
			r_v_2i_X_deg_chk_bit_b <= 0;
			
			r_EXECUTE_PE_DC <= 0;
	
			r_EXECUTE_PE_ELU <= 0;
			
			r_delta_2im2[`D_KES_GF_ORDER-1:0] <= D_KES_VALUE_ONE[`D_KES_GF_ORDER-1:0];
			
			r_delta_2im2_d0[`D_KES_GF_ORDER-1:0] <= 0;
		end
		
		else begin		
			case (r_nxt_state)
			KES_RESET: begin
				r_count_kes <= 0;
				r_sdr_buffer[(`D_KES_ECC_T*2*`D_KES_GF_ORDER)-1:0] <= 0;
				r_RESET_kes_sequence <= 1;
				
				r_v_2i_X_deg_chk_bit_b <= 0;
				
				r_EXECUTE_PE_DC <= 0;
		
				r_EXECUTE_PE_ELU <= 0;
				
				r_delta_2im2[`D_KES_GF_ORDER-1:0] <= D_KES_VALUE_ONE[`D_KES_GF_ORDER-1:0];
				
				r_delta_2im2_d0[`D_KES_GF_ORDER-1:0] <= 0;
			end
			KES_START: begin
				r_count_kes <= 0;
				/////////////////////////////////////////////
				////////// GENERATED BY C PROGRAMA //////////
				/////
				///
				
				// syndrome capture
					
				// buffer size: 1+63

				r_sdr_buffer[(`D_KES_ECC_T*2*`D_KES_GF_ORDER)-1:0] <= { D_KES_VALUE_ONE[`D_KES_GF_ORDER-1:0], i_syndromes[`D_KES_GF_ORDER*(`D_KES_ECC_T*2-1)-1:0] };

				                                          ///
														/////	
				////////// GENERATED BY C PROGRAMA //////////
				/////////////////////////////////////////////
				r_RESET_kes_sequence <= 0;
				
				r_v_2i_X_deg_chk_bit_b[`D_KES_ECC_T+1:0] <= w_v_2ip2_deg_info[`D_KES_ECC_T+1:0];
				
				r_EXECUTE_PE_DC <= 1;
		
				r_EXECUTE_PE_ELU <= 0;
				
				r_delta_2im2[`D_KES_GF_ORDER-1:0] <= w_delta_2i[`D_KES_GF_ORDER-1:0];
				
                r_delta_2im2_d0[`D_KES_GF_ORDER-1:0] <= 0;
			end
			KES_STEP1: begin
				r_count_kes <= r_count_kes + 1;
				r_sdr_buffer[(`D_KES_ECC_T*2*`D_KES_GF_ORDER)-1:0] <= r_sdr_buffer[(`D_KES_ECC_T*2*`D_KES_GF_ORDER)-1:0];
				r_RESET_kes_sequence <= 0;
				
				r_v_2i_X_deg_chk_bit_b[`D_KES_ECC_T+1:0] <= w_v_2ip2_deg_info[`D_KES_ECC_T+1:0];
				
				r_EXECUTE_PE_DC <= 0;
		
				r_EXECUTE_PE_ELU <= 1;
				
				r_delta_2im2[`D_KES_GF_ORDER-1:0] <= w_delta_2i[`D_KES_GF_ORDER-1:0];
				
				r_delta_2im2_d0[`D_KES_GF_ORDER-1:0] <= r_delta_2im2[`D_KES_GF_ORDER-1:0];
			end
			KES_STEP2: begin
				r_count_kes <= r_count_kes;
				r_sdr_buffer[(`D_KES_ECC_T*2*`D_KES_GF_ORDER)-1:0] <= (r_sdr_buffer[(`D_KES_ECC_T*2*`D_KES_GF_ORDER)-1:0]) << (`D_KES_GF_ORDER*2);
				r_RESET_kes_sequence <= 0;
				
				r_v_2i_X_deg_chk_bit_b[`D_KES_ECC_T+1:0] <= w_v_2ip2_deg_info[`D_KES_ECC_T+1:0];
				
				r_EXECUTE_PE_DC <= 1;
		
				r_EXECUTE_PE_ELU <= 0;
				
				r_delta_2im2[`D_KES_GF_ORDER-1:0] <= w_delta_2i[`D_KES_GF_ORDER-1:0];
				r_delta_2im2_d0 <= 0;
			end
            KES_FWD: begin
                r_count_kes <= 0;
				r_sdr_buffer[(`D_KES_ECC_T*2*`D_KES_GF_ORDER)-1:0] <= 0;
				r_RESET_kes_sequence <= 1;
				
				r_v_2i_X_deg_chk_bit_b <= 0;
				
				r_EXECUTE_PE_DC <= 0;
		
				r_EXECUTE_PE_ELU <= 0;
				
				r_delta_2im2[`D_KES_GF_ORDER-1:0] <= D_KES_VALUE_ONE[`D_KES_GF_ORDER-1:0];
				
				r_delta_2im2_d0[`D_KES_GF_ORDER-1:0] <= 0;
            end
            KES_PAUSE: begin
                r_count_kes <= r_count_kes;
				r_sdr_buffer[(`D_KES_ECC_T*2*`D_KES_GF_ORDER)-1:0] <= r_sdr_buffer[(`D_KES_ECC_T*2*`D_KES_GF_ORDER)-1:0];
				r_RESET_kes_sequence <= 0;
				
				r_v_2i_X_deg_chk_bit_b[`D_KES_ECC_T+1:0] <= r_v_2i_X_deg_chk_bit_b[`D_KES_ECC_T+1:0];
				
				r_EXECUTE_PE_DC <= 0;
		
				r_EXECUTE_PE_ELU <= 0;
				
				r_delta_2im2[`D_KES_GF_ORDER-1:0] <= r_delta_2im2[`D_KES_GF_ORDER-1:0];
				r_delta_2im2_d0 <= 0;
            end
			KES_OUT: begin
				r_count_kes <= r_count_kes;
				r_sdr_buffer[(`D_KES_ECC_T*2*`D_KES_GF_ORDER)-1:0] <= r_sdr_buffer[(`D_KES_ECC_T*2*`D_KES_GF_ORDER)-1:0];
				r_RESET_kes_sequence <= 0;
				
				r_v_2i_X_deg_chk_bit_b[`D_KES_ECC_T+1:0] <= r_v_2i_X_deg_chk_bit_b[`D_KES_ECC_T+1:0];
				
				r_EXECUTE_PE_DC <= 0;
		
				r_EXECUTE_PE_ELU <= 0;
				
				r_delta_2im2[`D_KES_GF_ORDER-1:0] <= r_delta_2im2[`D_KES_GF_ORDER-1:0];
				r_delta_2im2_d0 <= 0;
			end
			default: begin
				
			end
			endcase
		end
	end
	
	always @ (posedge i_clk)
	begin
		if ((i_RESET) || (i_stop_dec)) begin
            r_data_fowarding <= 0;
			o_chunk_number <= 0;
            o_channel_sel <= 0;
			o_buf_sequence_end <= 0;
			r_buf_sequence_end <= 0;
			end
		else begin
			case (r_nxt_state)
				KES_RESET: begin
                    r_data_fowarding <= 0;
					o_chunk_number <= 0;
                    o_channel_sel <= o_channel_sel;
					o_buf_sequence_end <= 0;
					r_buf_sequence_end <= 0;
					end
				KES_START: begin
                    r_data_fowarding <= i_data_fowarding;
					o_chunk_number <= i_chunk_number;
                    o_channel_sel <= i_channel_sel;
					o_buf_sequence_end <= 0;
					r_buf_sequence_end <= i_buf_sequence_end;
					end
				KES_OUT: begin
                    r_data_fowarding <= r_data_fowarding;
					o_chunk_number <= o_chunk_number;
                    o_channel_sel <= o_channel_sel;
					o_buf_sequence_end <= r_buf_sequence_end;
					r_buf_sequence_end <= r_buf_sequence_end;
					end
				default: begin
                    r_data_fowarding <= r_data_fowarding;
					o_chunk_number <= o_chunk_number;
                    o_channel_sel <= o_channel_sel;
					o_buf_sequence_end <= 0;
					r_buf_sequence_end <= r_buf_sequence_end;
					end
			endcase
			end
	end
	
	always @ (posedge i_clk)
	begin
		if ((i_RESET) || (i_stop_dec)) begin
			o_error_count <= 0;
			end
		else
			case (r_nxt_state)
				KES_OUT: begin
					casez (w_v_error[`D_KES_ECC_T:0])
						15'b1?????????????1: begin
							o_error_count <= 4'b1110;
						end
						15'b1????????????10: begin
							o_error_count <= 4'b1101;
						end
						15'b1???????????100: begin
							o_error_count <= 4'b1100;
						end
						15'b1??????????1000: begin
							o_error_count <= 4'b1011;
						end
						15'b1?????????10000: begin
							o_error_count <= 4'b1010;
						end
						15'b1????????100000: begin
							o_error_count <= 4'b1001;
						end
						15'b1???????1000000: begin
							o_error_count <= 4'b1000;
						end
						15'b1??????10000000: begin
							o_error_count <= 4'b0111;
						end
						15'b1?????100000000: begin
							o_error_count <= 4'b0110;
						end
						15'b1????1000000000: begin
							o_error_count <= 4'b0101;
						end
						15'b1???10000000000: begin
							o_error_count <= 4'b0100;
						end
						15'b1??100000000000: begin
							o_error_count <= 4'b0011;
						end
						15'b1?1000000000000: begin
							o_error_count <= 4'b0010;
						end
						15'b110000000000000: begin
							o_error_count <= 4'b0001;
						end
						default: begin
							o_error_count <= 4'b0000;
						end
						endcase
					end
			default:
				o_error_count <= 0;
			endcase
	end
	
	// MAXIMUM degree checker
	always @ (posedge i_clk)
	begin
		if ((w_RESET_KES) || (i_stop_dec)) begin
			r_ELP_degree_condition_violation <= 0;
			r_v_2i_maximum_deg[`D_KES_ECC_T_BIT-1:0] <= 0;
		end	else begin			
			/////////////////////////////////////////////
			////////// GENERATED BY C PROGRAMA //////////
			/////
			///
			
			// check maximum degree
			
			// violation check
			// casez: 34
			
			r_ELP_degree_condition_violation <= (w_last_interation)? r_v_2i_X_deg_chk_bit_b[`D_KES_ECC_T+1]:1'b0;

            casez (r_v_2i_X_deg_chk_bit_b[`D_KES_ECC_T+1:0])
            16'b000000000000000?: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b0000;
            end

            16'b000000000000001?: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b0001;
            end

            16'b00000000000001??: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b0010;
            end

            16'b0000000000001???: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b0011;
            end

            16'b000000000001????: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b0100;
            end

            16'b00000000001?????: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b0101;
            end

            16'b0000000001??????: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b0110;
            end

            16'b000000001???????: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b0111;
            end

            16'b00000001????????: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b1000;
            end

            16'b0000001?????????: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b1001;
            end

            16'b000001??????????: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b1010;
            end

            16'b00001???????????: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b1011;
            end

            16'b0001????????????: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b1100;
            end

            16'b001?????????????: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b1101;
            end

            16'b01??????????????: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b1110;
            end

            16'b1???????????????: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b1111;
            end
            default: begin
                r_v_2i_maximum_deg[`D_KES_ECC_T_BIT - 1:0] <= 4'b0000;
            end
            endcase
			
			                                          ///
													/////	
			////////// GENERATED BY C PROGRAMA //////////
			/////////////////////////////////////////////
		end
	end
	
	
	
	// processing elements
	
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// PE_DC, PE_ELU
	
	// sdr_connection_wire: 31, t+1-2
	// PE_DC: 33, t+1
	// k: 33 t+2-1
	// PE_ELU: 34, t+2
	
    
    wire [`D_KES_GF_ORDER-1:0] w_sdr_from_DC_012_to_DC_014;
    wire [`D_KES_GF_ORDER-1:0] w_sdr_from_DC_011_to_DC_013;
    wire [`D_KES_GF_ORDER-1:0] w_sdr_from_DC_010_to_DC_012;
    wire [`D_KES_GF_ORDER-1:0] w_sdr_from_DC_009_to_DC_011;
    wire [`D_KES_GF_ORDER-1:0] w_sdr_from_DC_008_to_DC_010;
    wire [`D_KES_GF_ORDER-1:0] w_sdr_from_DC_007_to_DC_009;
    wire [`D_KES_GF_ORDER-1:0] w_sdr_from_DC_006_to_DC_008;
    wire [`D_KES_GF_ORDER-1:0] w_sdr_from_DC_005_to_DC_007;
    wire [`D_KES_GF_ORDER-1:0] w_sdr_from_DC_004_to_DC_006;
    wire [`D_KES_GF_ORDER-1:0] w_sdr_from_DC_003_to_DC_005;
    wire [`D_KES_GF_ORDER-1:0] w_sdr_from_DC_002_to_DC_004;
    wire [`D_KES_GF_ORDER-1:0] w_sdr_from_DC_001_to_DC_003;
    wire [`D_KES_GF_ORDER-1:0] w_sdr_from_DC_000_to_DC_002;

    d_KES_PE_DC_2MAXodr DC_014 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_from_DC_012_to_DC_014[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_014[`D_KES_GF_ORDER-1:0]),

    .o_coef_2ip1(w_coef_2ip1_014[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_2MAXodr DC_013 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_from_DC_011_to_DC_013[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_013[`D_KES_GF_ORDER-1:0]),

    .o_coef_2ip1(w_coef_2ip1_013[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_NMLodr DC_012 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_from_DC_010_to_DC_012[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_012[`D_KES_GF_ORDER-1:0]),

    .o_S_out(w_sdr_from_DC_012_to_DC_014[`D_KES_GF_ORDER - 1:0]),
    .o_coef_2ip1(w_coef_2ip1_012[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_NMLodr DC_011 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_from_DC_009_to_DC_011[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_011[`D_KES_GF_ORDER-1:0]),

    .o_S_out(w_sdr_from_DC_011_to_DC_013[`D_KES_GF_ORDER - 1:0]),
    .o_coef_2ip1(w_coef_2ip1_011[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_NMLodr DC_010 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_from_DC_008_to_DC_010[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_010[`D_KES_GF_ORDER-1:0]),

    .o_S_out(w_sdr_from_DC_010_to_DC_012[`D_KES_GF_ORDER - 1:0]),
    .o_coef_2ip1(w_coef_2ip1_010[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_NMLodr DC_009 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_from_DC_007_to_DC_009[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_009[`D_KES_GF_ORDER-1:0]),

    .o_S_out(w_sdr_from_DC_009_to_DC_011[`D_KES_GF_ORDER - 1:0]),
    .o_coef_2ip1(w_coef_2ip1_009[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_NMLodr DC_008 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_from_DC_006_to_DC_008[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_008[`D_KES_GF_ORDER-1:0]),

    .o_S_out(w_sdr_from_DC_008_to_DC_010[`D_KES_GF_ORDER - 1:0]),
    .o_coef_2ip1(w_coef_2ip1_008[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_NMLodr DC_007 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_from_DC_005_to_DC_007[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_007[`D_KES_GF_ORDER-1:0]),

    .o_S_out(w_sdr_from_DC_007_to_DC_009[`D_KES_GF_ORDER - 1:0]),
    .o_coef_2ip1(w_coef_2ip1_007[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_NMLodr DC_006 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_from_DC_004_to_DC_006[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_006[`D_KES_GF_ORDER-1:0]),

    .o_S_out(w_sdr_from_DC_006_to_DC_008[`D_KES_GF_ORDER - 1:0]),
    .o_coef_2ip1(w_coef_2ip1_006[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_NMLodr DC_005 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_from_DC_003_to_DC_005[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_005[`D_KES_GF_ORDER-1:0]),

    .o_S_out(w_sdr_from_DC_005_to_DC_007[`D_KES_GF_ORDER - 1:0]),
    .o_coef_2ip1(w_coef_2ip1_005[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_NMLodr DC_004 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_from_DC_002_to_DC_004[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_004[`D_KES_GF_ORDER-1:0]),

    .o_S_out(w_sdr_from_DC_004_to_DC_006[`D_KES_GF_ORDER - 1:0]),
    .o_coef_2ip1(w_coef_2ip1_004[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_NMLodr DC_003 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_from_DC_001_to_DC_003[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_003[`D_KES_GF_ORDER-1:0]),

    .o_S_out(w_sdr_from_DC_003_to_DC_005[`D_KES_GF_ORDER - 1:0]),
    .o_coef_2ip1(w_coef_2ip1_003[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_NMLodr DC_002 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_from_DC_000_to_DC_002[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_002[`D_KES_GF_ORDER-1:0]),

    .o_S_out(w_sdr_from_DC_002_to_DC_004[`D_KES_GF_ORDER - 1:0]),
    .o_coef_2ip1(w_coef_2ip1_002[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_NMLodr DC_001 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_to_DC_001[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_001[`D_KES_GF_ORDER-1:0]),

    .o_S_out(w_sdr_from_DC_001_to_DC_003[`D_KES_GF_ORDER - 1:0]),
    .o_coef_2ip1(w_coef_2ip1_001[`D_KES_GF_ORDER - 1:0]));

    d_KES_PE_DC_NMLodr DC_000 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
	.i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_DC(r_EXECUTE_PE_DC),
    .i_S_in(w_sdr_to_DC_000[`D_KES_GF_ORDER - 1:0]),
    .i_v_2i_X(o_v_2i_000[`D_KES_GF_ORDER-1:0]),

    .o_S_out(w_sdr_from_DC_000_to_DC_002[`D_KES_GF_ORDER - 1:0]),
    .o_coef_2ip1(w_coef_2ip1_000[`D_KES_GF_ORDER - 1:0]));
	
   
    
    wire [`D_KES_GF_ORDER-1:0] w_k_014;
    wire [`D_KES_GF_ORDER-1:0] w_k_013;
    wire [`D_KES_GF_ORDER-1:0] w_k_012;
    wire [`D_KES_GF_ORDER-1:0] w_k_011;
    wire [`D_KES_GF_ORDER-1:0] w_k_010;
    wire [`D_KES_GF_ORDER-1:0] w_k_009;
    wire [`D_KES_GF_ORDER-1:0] w_k_008;
    wire [`D_KES_GF_ORDER-1:0] w_k_007;
    wire [`D_KES_GF_ORDER-1:0] w_k_006;
    wire [`D_KES_GF_ORDER-1:0] w_k_005;
    wire [`D_KES_GF_ORDER-1:0] w_k_004;
    wire [`D_KES_GF_ORDER-1:0] w_k_003;
    wire [`D_KES_GF_ORDER-1:0] w_k_002;
    wire [`D_KES_GF_ORDER-1:0] w_k_001;
    wire [`D_KES_GF_ORDER-1:0] w_k_000;

    d_KES_PE_ELU_eMAXodr ELU_015 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_k_2i_Xm1(w_k_014[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),

    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_015));

    d_KES_PE_ELU_NMLodr ELU_014 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_013[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_013[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm2(w_k_012[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_014[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_014),
    .o_k_2i_X(w_k_014[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_NMLodr ELU_013 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_012[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_012[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm2(w_k_011[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_013[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_013),
    .o_k_2i_X(w_k_013[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_NMLodr ELU_012 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_011[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_011[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm2(w_k_010[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_012[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_012),
    .o_k_2i_X(w_k_012[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_NMLodr ELU_011 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_010[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_010[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm2(w_k_009[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_011[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_011),
    .o_k_2i_X(w_k_011[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_NMLodr ELU_010 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_009[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_009[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm2(w_k_008[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_010[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_010),
    .o_k_2i_X(w_k_010[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_NMLodr ELU_009 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_008[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_008[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm2(w_k_007[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_009[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_009),
    .o_k_2i_X(w_k_009[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_NMLodr ELU_008 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_007[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_007[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm2(w_k_006[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_008[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_008),
    .o_k_2i_X(w_k_008[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_NMLodr ELU_007 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_006[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_006[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm2(w_k_005[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_007[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_007),
    .o_k_2i_X(w_k_007[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_NMLodr ELU_006 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_005[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_005[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm2(w_k_004[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_006[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_006),
    .o_k_2i_X(w_k_006[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_NMLodr ELU_005 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_004[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_004[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm2(w_k_003[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_005[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_005),
    .o_k_2i_X(w_k_005[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_NMLodr ELU_004 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_003[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_003[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm2(w_k_002[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_004[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_004),
    .o_k_2i_X(w_k_004[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_NMLodr ELU_003 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_002[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_002[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm2(w_k_001[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_003[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_003),
    .o_k_2i_X(w_k_003[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_NMLodr ELU_002 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_001[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_001[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm2(w_k_000[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_002[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_002),
    .o_k_2i_X(w_k_002[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_sMINodr ELU_001 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_v_2i_Xm1(o_v_2i_000[`D_KES_GF_ORDER-1:0]),
    .i_k_2i_Xm1(w_k_000[`D_KES_GF_ORDER-1:0]),
    .i_d_2i(w_d_2i[`D_KES_GF_ORDER-1:0]),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),
    .i_condition_2i(w_condition_2i),

    .o_v_2i_X(o_v_2i_001[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_001),
    .o_k_2i_X(w_k_001[`D_KES_GF_ORDER-1:0]));

    d_KES_PE_ELU_MINodr ELU_000 (
    .i_clk(i_clk),
    .i_RESET_KES(w_RESET_KES),
    .i_stop_dec(i_stop_dec),
    .i_EXECUTE_PE_ELU(r_EXECUTE_PE_ELU),
    .i_delta_2im2(r_delta_2im2_d0[`D_KES_GF_ORDER-1:0]),

    .o_v_2i_X(o_v_2i_000[`D_KES_GF_ORDER-1:0]),
    .o_v_2i_X_deg_chk_bit(w_v_2i_X_deg_chk_bit_000),
    .o_k_2i_X(w_k_000[`D_KES_GF_ORDER-1:0]));
	
	                                          ///
											/////	
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
	
	
endmodule
