

`include "d_CS_parameters.vh"
`timescale 1ns / 1ps

module d_BCH_CS_top
(
	input  wire                       i_clk,
    input  wire                       i_RESET,
    input  wire						  i_stop_dec,
	
	output wire                       o_cs_available,           // [indicate] Chien search ready
	
	input  wire                       i_exe_cs,                 // Chien search start command signal
    input  wire                       i_data_fowarding,        
	input  wire						  i_MUX_data_ready,				
	
	
	output wire                       o_cs_start,               // [indicate] Chien search start
	output wire                       o_cs_cmplt,               // [indicate] Chien search complete
	output wire						  o_cs_pause,				// [indicate] Ch
	
	output wire                       o_BRAM_read_enable,
	output wire [`D_CS_O_CNT_BIT-2:0] o_BRAM_read_address,
	input  wire [`D_CS_P_LVL-1:0]     i_BRAM_read_data,         // received code
	
	output wire                       o_c_message_valid,        // [indicate] corrected message BUS strobe signal
    output wire                       o_c_message_output_start, // [indicate] corrected message output start
    output wire                       o_c_message_output_cmplt, // [indicate] corrected message output complete
	
    output reg  [`D_CS_P_LVL-1:0]     o_c_message,              // corrected message BUS
	
	
	
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// total: 15
	
	input wire [`D_CS_GF_ORDER-1:0] i_v_000,
    input wire [`D_CS_GF_ORDER-1:0] i_v_001,
    input wire [`D_CS_GF_ORDER-1:0] i_v_002,
    input wire [`D_CS_GF_ORDER-1:0] i_v_003,
    input wire [`D_CS_GF_ORDER-1:0] i_v_004,
    input wire [`D_CS_GF_ORDER-1:0] i_v_005,
    input wire [`D_CS_GF_ORDER-1:0] i_v_006,
    input wire [`D_CS_GF_ORDER-1:0] i_v_007,
    input wire [`D_CS_GF_ORDER-1:0] i_v_008,
    input wire [`D_CS_GF_ORDER-1:0] i_v_009,
    input wire [`D_CS_GF_ORDER-1:0] i_v_010,
    input wire [`D_CS_GF_ORDER-1:0] i_v_011,
    input wire [`D_CS_GF_ORDER-1:0] i_v_012,
    input wire [`D_CS_GF_ORDER-1:0] i_v_013,
    input wire [`D_CS_GF_ORDER-1:0] i_v_014
    
	
	                                          ///
	                                        /////
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
    );
	
	parameter CS_FSM_BIT = 13;
	parameter RESET      = 13'b0000000000001; // RESET
    parameter DELAY      = 13'b0000000000010;
    parameter DELAY_FWD  = 13'b0000000000100;
	parameter EVAL_SHT   = 13'b0000000001000; // evaluation shortening
	parameter CS_STRT    = 13'b0000000010000; // Chien search, start
	parameter CS_FBCK    = 13'b0000000100000; // Chien search, feedback
	parameter CS_STBY	 = 13'b0000001000000; // Chien search, pause
	parameter CS_FNLS    = 13'b0000010000000; // final stage, output last corrected message
    parameter FWD_MODE   = 13'b0000100000000;
    parameter FWD_STRT   = 13'b0001000000000; // Forwarding, Correction is not needed or possible
    parameter FWD_FBCK   = 13'b0010000000000; // Forwarding
    parameter FWD_STBY   = 13'b0100000000000; // Forwarding
    parameter FWD_FNLS   = 13'b1000000000000; // Forwarding
	
	
	
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// total: 8, 8
	
	wire w_slot_001_flip;
    wire w_slot_002_flip;
    wire w_slot_003_flip;
    wire w_slot_004_flip;
    wire w_slot_005_flip;
    wire w_slot_006_flip;
    wire w_slot_007_flip;
    wire w_slot_008_flip;

    wire w_slot_001_flipped_message;
    wire w_slot_002_flipped_message;
    wire w_slot_003_flipped_message;
    wire w_slot_004_flipped_message;
    wire w_slot_005_flipped_message;
    wire w_slot_006_flipped_message;
    wire w_slot_007_flipped_message;
    wire w_slot_008_flipped_message;
	
	                                          ///
	                                        /////
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
	
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// total: 14
	
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_001;
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_002;
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_003;
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_004;
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_005;
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_006;
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_007;
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_008;
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_009;
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_010;
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_011;
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_012;
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_013;
    wire [`D_CS_GF_ORDER -1:0] w_shortened_v_014;
	
	                                          ///
	                                        /////
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
	
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// total: 15
	
	wire [`D_CS_GF_ORDER -1:0] w_ELP_term_000;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_001;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_002;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_003;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_004;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_005;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_006;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_007;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_008;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_009;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_010;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_011;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_012;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_013;
    wire [`D_CS_GF_ORDER -1:0] w_ELP_term_014;
	
	                                          ///
	                                        /////
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
	
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// total: 15 * 8 = 120
	
	wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_000;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_001;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_002;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_003;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_004;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_005;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_006;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_007;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_008;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_009;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_010;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_011;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_012;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_013;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S001_014;

    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_000;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_001;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_002;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_003;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_004;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_005;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_006;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_007;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_008;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_009;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_010;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_011;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_012;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_013;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S002_014;

    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_000;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_001;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_002;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_003;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_004;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_005;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_006;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_007;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_008;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_009;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_010;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_011;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_012;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_013;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S003_014;

    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_000;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_001;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_002;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_003;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_004;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_005;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_006;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_007;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_008;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_009;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_010;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_011;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_012;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_013;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S004_014;

    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_000;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_001;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_002;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_003;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_004;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_005;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_006;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_007;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_008;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_009;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_010;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_011;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_012;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_013;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S005_014;

    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_000;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_001;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_002;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_003;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_004;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_005;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_006;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_007;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_008;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_009;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_010;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_011;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_012;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_013;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S006_014;

    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_000;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_001;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_002;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_003;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_004;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_005;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_006;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_007;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_008;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_009;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_010;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_011;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_012;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_013;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S007_014;

    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_000;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_001;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_002;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_003;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_004;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_005;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_006;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_007;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_008;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_009;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_010;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_011;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_012;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_013;
    wire [`D_CS_GF_ORDER-1:0] w_evaluated_term_S008_014;
    
	
	                                          ///
	                                        /////
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
	
	// encoder FSM state
	reg  [CS_FSM_BIT-1:0] r_cur_state;
	reg  [CS_FSM_BIT-1:0] r_nxt_state;
	
	// internal counter
	reg  [`D_CS_O_CNT_BIT:0] r_counter;
	
	// internal variable
	wire [(`D_CS_ECC_T+1)*`D_CS_GF_ORDER -1:`D_CS_GF_ORDER ] w_v_input_wire_e000; // i_v_014 ~ i_v_001, except i_v_000
	reg  [(`D_CS_ECC_T+1)*`D_CS_GF_ORDER -1:`D_CS_GF_ORDER ] r_v_buffer_e000;     // i_v_014 ~ i_v_001, except i_v_000
    reg  [(`D_CS_ECC_T+1)*`D_CS_GF_ORDER -1:`D_CS_GF_ORDER ] r_v_buffer_e000_delay;  

    
	reg  [`D_CS_GF_ORDER -1:0]                               r_v_buffer_000;      // i_v_000
    reg  [`D_CS_GF_ORDER -1:0]                               r_v_buffer_000_delay;
	
	wire [(`D_CS_ECC_T+1)*`D_CS_GF_ORDER -1:`D_CS_GF_ORDER ] w_shortened_v;       // i_v_014 ~ i_v_001
	wire [(`D_CS_ECC_T+1)*`D_CS_GF_ORDER -1:`D_CS_GF_ORDER ] w_feedback_wire;     // i_v_014 ~ i_v_001
	
	reg  [(`D_CS_ECC_T+1)*`D_CS_GF_ORDER -1:`D_CS_GF_ORDER ] r_feedback_buffer;   // i_v_014 ~ i_v_001
	
	reg  [`D_CS_P_LVL-1:0] r_received_code_buffer;
    reg  [`D_CS_P_LVL-1:0] r_BRAM_read_buffer;
    reg  [`D_CS_P_LVL-1:0] r_waiting_buffer;
	wire [`D_CS_P_LVL-1:0] w_flipped_message;
	
	
	
	// generate control/indicate signal
	assign o_BRAM_read_enable = (i_exe_cs) | ( ((r_cur_state == DELAY) | (r_cur_state == DELAY_FWD) | (r_cur_state == EVAL_SHT) | (r_cur_state == CS_STRT) | (r_cur_state == CS_FBCK) | (r_cur_state == FWD_MODE) | (r_cur_state == FWD_STRT) | (r_cur_state == FWD_FBCK)) & (r_counter != `D_CS_O_CNT) & (r_counter != `D_CS_O_CNT+1) & (r_counter != `D_CS_O_CNT+2) );
	assign o_BRAM_read_address = r_counter[`D_CS_O_CNT_BIT-2:0];
	
	assign o_cs_start = (r_cur_state == EVAL_SHT) || (r_cur_state == FWD_MODE);
	assign o_cs_available = (r_cur_state == RESET);
	assign o_cs_cmplt = ((r_cur_state == CS_FNLS) | (r_cur_state == FWD_FNLS)) & i_MUX_data_ready & o_c_message_valid;
	
	assign o_c_message_valid = (r_cur_state == CS_FBCK) | (r_cur_state == CS_FNLS) | (r_cur_state == CS_STBY) | (r_cur_state == FWD_FBCK) | (r_cur_state == FWD_FNLS) | (r_cur_state == FWD_STBY) ;
	assign o_c_message_output_start = (r_counter == 4);
	assign o_c_message_output_cmplt = o_cs_cmplt;
	assign o_cs_pause = (r_cur_state == CS_STBY) || (r_cur_state == FWD_STBY);

	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// wire mapping
	
	assign w_v_input_wire_e000[(`D_CS_ECC_T+1)*`D_CS_GF_ORDER-1:`D_CS_GF_ORDER] = { i_v_014[`D_CS_GF_ORDER-1:0], i_v_013[`D_CS_GF_ORDER-1:0], i_v_012[`D_CS_GF_ORDER-1:0], i_v_011[`D_CS_GF_ORDER-1:0], i_v_010[`D_CS_GF_ORDER-1:0], i_v_009[`D_CS_GF_ORDER-1:0], i_v_008[`D_CS_GF_ORDER-1:0], i_v_007[`D_CS_GF_ORDER-1:0], i_v_006[`D_CS_GF_ORDER-1:0], i_v_005[`D_CS_GF_ORDER-1:0], i_v_004[`D_CS_GF_ORDER-1:0], i_v_003[`D_CS_GF_ORDER-1:0], i_v_002[`D_CS_GF_ORDER-1:0], i_v_001[`D_CS_GF_ORDER-1:0] };

    assign w_shortened_v[(`D_CS_ECC_T+1)*`D_CS_GF_ORDER-1:`D_CS_GF_ORDER] = { w_shortened_v_014[`D_CS_GF_ORDER-1:0], w_shortened_v_013[`D_CS_GF_ORDER-1:0], w_shortened_v_012[`D_CS_GF_ORDER-1:0], w_shortened_v_011[`D_CS_GF_ORDER-1:0], w_shortened_v_010[`D_CS_GF_ORDER-1:0], w_shortened_v_009[`D_CS_GF_ORDER-1:0], w_shortened_v_008[`D_CS_GF_ORDER-1:0], w_shortened_v_007[`D_CS_GF_ORDER-1:0], w_shortened_v_006[`D_CS_GF_ORDER-1:0], w_shortened_v_005[`D_CS_GF_ORDER-1:0], w_shortened_v_004[`D_CS_GF_ORDER-1:0], w_shortened_v_003[`D_CS_GF_ORDER-1:0], w_shortened_v_002[`D_CS_GF_ORDER-1:0], w_shortened_v_001[`D_CS_GF_ORDER-1:0] };

    assign w_feedback_wire[(`D_CS_ECC_T+1)*`D_CS_GF_ORDER-1:`D_CS_GF_ORDER] = { w_evaluated_term_S008_014[`D_CS_GF_ORDER-1:0], w_evaluated_term_S008_013[`D_CS_GF_ORDER-1:0], w_evaluated_term_S008_012[`D_CS_GF_ORDER-1:0], w_evaluated_term_S008_011[`D_CS_GF_ORDER-1:0], w_evaluated_term_S008_010[`D_CS_GF_ORDER-1:0], w_evaluated_term_S008_009[`D_CS_GF_ORDER-1:0], w_evaluated_term_S008_008[`D_CS_GF_ORDER-1:0], w_evaluated_term_S008_007[`D_CS_GF_ORDER-1:0], w_evaluated_term_S008_006[`D_CS_GF_ORDER-1:0], w_evaluated_term_S008_005[`D_CS_GF_ORDER-1:0], w_evaluated_term_S008_004[`D_CS_GF_ORDER-1:0], w_evaluated_term_S008_003[`D_CS_GF_ORDER-1:0], w_evaluated_term_S008_002[`D_CS_GF_ORDER-1:0], w_evaluated_term_S008_001[`D_CS_GF_ORDER-1:0] };

	                                          ///
	                                        /////
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
	
	assign w_ELP_term_000[`D_CS_GF_ORDER -1:0] = r_v_buffer_000[`D_CS_GF_ORDER -1:0];
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// total: 14
	
    
	assign w_ELP_term_001[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[(  1+1)*`D_CS_GF_ORDER-1:(  1+0)*`D_CS_GF_ORDER];
    assign w_ELP_term_002[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[(  2+1)*`D_CS_GF_ORDER-1:(  2+0)*`D_CS_GF_ORDER];
    assign w_ELP_term_003[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[(  3+1)*`D_CS_GF_ORDER-1:(  3+0)*`D_CS_GF_ORDER];
    assign w_ELP_term_004[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[(  4+1)*`D_CS_GF_ORDER-1:(  4+0)*`D_CS_GF_ORDER];
    assign w_ELP_term_005[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[(  5+1)*`D_CS_GF_ORDER-1:(  5+0)*`D_CS_GF_ORDER];
    assign w_ELP_term_006[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[(  6+1)*`D_CS_GF_ORDER-1:(  6+0)*`D_CS_GF_ORDER];
    assign w_ELP_term_007[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[(  7+1)*`D_CS_GF_ORDER-1:(  7+0)*`D_CS_GF_ORDER];
    assign w_ELP_term_008[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[(  8+1)*`D_CS_GF_ORDER-1:(  8+0)*`D_CS_GF_ORDER];
    assign w_ELP_term_009[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[(  9+1)*`D_CS_GF_ORDER-1:(  9+0)*`D_CS_GF_ORDER];
    assign w_ELP_term_010[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[( 10+1)*`D_CS_GF_ORDER-1:( 10+0)*`D_CS_GF_ORDER];
    assign w_ELP_term_011[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[( 11+1)*`D_CS_GF_ORDER-1:( 11+0)*`D_CS_GF_ORDER];
    assign w_ELP_term_012[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[( 12+1)*`D_CS_GF_ORDER-1:( 12+0)*`D_CS_GF_ORDER];
    assign w_ELP_term_013[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[( 13+1)*`D_CS_GF_ORDER-1:( 13+0)*`D_CS_GF_ORDER];
    assign w_ELP_term_014[`D_CS_GF_ORDER-1:0] = r_feedback_buffer[( 14+1)*`D_CS_GF_ORDER-1:( 14+0)*`D_CS_GF_ORDER];
	
	                                          ///
	                                        /////
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
	
	
		
	// update current state to next state
	always @ (posedge i_clk)
	begin
		if ((i_RESET) || (i_stop_dec))
			r_cur_state <= RESET;
		else
			r_cur_state <= r_nxt_state;
	end
	
	// decide next state
	always @ ( * )
	begin
		case (r_cur_state)
		RESET: begin
			r_nxt_state <= (i_exe_cs)? ((i_data_fowarding)? DELAY_FWD:DELAY):RESET;
		end
        DELAY: begin
            r_nxt_state <= EVAL_SHT;
        end
		EVAL_SHT: begin
			r_nxt_state <= CS_STRT;
		end
		CS_STRT: begin
			r_nxt_state <= CS_FBCK;
		end
		CS_FBCK: begin
			r_nxt_state <= (!i_MUX_data_ready)? CS_STBY : ((r_counter == `D_CS_O_CNT+2)? (CS_FNLS):(CS_FBCK));
		end
		CS_STBY:	begin
			r_nxt_state <= (!i_MUX_data_ready)? CS_STBY: ((r_counter == `D_CS_O_CNT+2)? CS_FNLS: CS_FBCK);
		end
		CS_FNLS: begin
			r_nxt_state <= (!i_MUX_data_ready)? CS_FNLS: ((i_exe_cs)? ((i_data_fowarding)? FWD_MODE:EVAL_SHT):RESET);
		end
        DELAY_FWD: begin
            r_nxt_state <= FWD_MODE;
        end
        FWD_MODE: begin
            r_nxt_state <= FWD_STRT;
        end
        FWD_STRT: begin
            r_nxt_state <= FWD_FBCK;
        end
        FWD_FBCK: begin
            r_nxt_state <= (!i_MUX_data_ready)? FWD_STBY : ((r_counter == `D_CS_O_CNT+2)? (FWD_FNLS):(FWD_FBCK));
        end
        FWD_STBY: begin
            r_nxt_state <= (!i_MUX_data_ready)? FWD_STBY : ((r_counter == `D_CS_O_CNT+2)? (FWD_FNLS):(FWD_FBCK));
        end
        FWD_FNLS: begin
            r_nxt_state <= (!i_MUX_data_ready)? FWD_FNLS : ((i_exe_cs)? ((i_data_fowarding)? FWD_MODE:EVAL_SHT):RESET);
        end
		default: begin
			r_nxt_state <= RESET;
		end
		endcase
	end
	
	// state behaviour
	always @ (posedge i_clk)
	begin
			case (r_nxt_state)
			
			RESET:begin
				r_counter <= 0;
				
                r_v_buffer_e000_delay <= 0;
                r_v_buffer_000_delay <= 0;
                
				r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= 0;
				
				r_feedback_buffer <= 0;
				
                r_BRAM_read_buffer <= 0;
                r_waiting_buffer <= 0;
				r_received_code_buffer <= 0;
				o_c_message <= 0;
			end
			
            DELAY: begin
                r_counter <= 1;
                
                r_v_buffer_e000_delay <= w_v_input_wire_e000;
                r_v_buffer_000_delay <= i_v_000;
                
                r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= 0;
				
				r_feedback_buffer <= 0;
				
                r_BRAM_read_buffer <= 0;
                r_waiting_buffer <= 0;
				r_received_code_buffer <= 0;
				o_c_message <= 0;
            end
            
			EVAL_SHT: begin
				r_counter <= 2;
				
                r_v_buffer_e000_delay <= 0;
                r_v_buffer_000_delay <= r_v_buffer_000_delay;
                
				r_v_buffer_e000 <= r_v_buffer_e000_delay;
				r_v_buffer_000 <= r_v_buffer_000_delay;
				
				r_feedback_buffer <= 0;
				
                r_BRAM_read_buffer <= i_BRAM_read_data;
                r_waiting_buffer <= i_BRAM_read_data;
				r_received_code_buffer <= 0;
				o_c_message <= 0;
			end
			
			CS_STRT: begin
				r_counter <= 3;
				
                r_v_buffer_e000_delay <= 0;
                r_v_buffer_000_delay <= 0;
                
				r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= r_v_buffer_000;
				
				r_feedback_buffer <= w_shortened_v;
				
                r_BRAM_read_buffer <= i_BRAM_read_data;
                r_waiting_buffer <= i_BRAM_read_data;
				r_received_code_buffer <= r_BRAM_read_buffer;
				o_c_message <= 0;
			end
			
			CS_FBCK:
            begin
                r_counter <= r_counter + 1'b1;
				
                r_v_buffer_e000_delay <= 0;
                r_v_buffer_000_delay <= 0;
                
				r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= r_v_buffer_000;
				
				r_feedback_buffer <= w_feedback_wire;
				
                r_BRAM_read_buffer <= i_BRAM_read_data;
                r_waiting_buffer <= (r_cur_state == CS_STBY) ? r_BRAM_read_buffer:i_BRAM_read_data;
				r_received_code_buffer <= r_waiting_buffer;
				o_c_message <= w_flipped_message;
            end
                
			
			
			CS_STBY:
            begin
                r_counter <= r_counter;
				
                r_v_buffer_e000_delay <= 0;
                r_v_buffer_000_delay <= 0;
                
				r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= r_v_buffer_000;
				
				r_feedback_buffer <= r_feedback_buffer;
				
                r_BRAM_read_buffer <= (r_cur_state == CS_STBY)? r_BRAM_read_buffer:i_BRAM_read_data;
                r_waiting_buffer <= r_waiting_buffer;
				r_received_code_buffer <= r_received_code_buffer;
                
				o_c_message <= o_c_message;
            end
			
			CS_FNLS: begin
			if (r_cur_state == CS_FNLS) begin
				r_counter <= 0;
				
				r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= 0;
				
				r_feedback_buffer <= 0;
				
				r_received_code_buffer <= 0;
				o_c_message <= o_c_message;
				end
			else begin
				r_counter <= 0;
				
				r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= 0;
				
				r_feedback_buffer <= 0;
				
				r_received_code_buffer <= 0;
				o_c_message <= w_flipped_message;
				end
			end
            DELAY_FWD: begin
                r_counter <= 1;
                
                r_v_buffer_e000_delay <= w_v_input_wire_e000;
                r_v_buffer_000_delay <= i_v_000;
                
                r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= 0;
				
				r_feedback_buffer <= 0;
				
                r_BRAM_read_buffer <= 0;
                r_waiting_buffer <= 0;
				r_received_code_buffer <= 0;
				o_c_message <= 0;
            end
            FWD_MODE: begin
				r_counter <= 2;
				
                r_v_buffer_e000_delay <= 0;
                r_v_buffer_000_delay <= r_v_buffer_000_delay;
                
				r_v_buffer_e000 <= r_v_buffer_e000_delay;
				r_v_buffer_000 <= r_v_buffer_000_delay;
				
				r_feedback_buffer <= 0;
				
                r_BRAM_read_buffer <= i_BRAM_read_data;
                r_waiting_buffer <= i_BRAM_read_data;
				r_received_code_buffer <= 0;
				o_c_message <= 0;
			end
            
			FWD_STRT: begin
                r_counter <= 3;
				
                r_v_buffer_e000_delay <= 0;
                r_v_buffer_000_delay <= 0;
                
				r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= 0;
				
				r_feedback_buffer <= 0;
				
                r_BRAM_read_buffer <= i_BRAM_read_data;
                r_waiting_buffer <= i_BRAM_read_data;
				r_received_code_buffer <= r_BRAM_read_buffer;
				o_c_message <= 0;
			end
            
            FWD_FBCK: begin
				r_counter <= r_counter + 1'b1;
				
				r_v_buffer_e000_delay <= 0;
                r_v_buffer_000_delay <= 0;
                
				r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= 0;
				
				r_feedback_buffer <= 0;
				
                r_BRAM_read_buffer <= i_BRAM_read_data;
                r_waiting_buffer <= (r_cur_state == FWD_STBY) ? r_BRAM_read_buffer:i_BRAM_read_data;
				r_received_code_buffer <= r_waiting_buffer;
				o_c_message <= r_received_code_buffer;
			end
            FWD_STBY: begin
				r_counter <= r_counter;
				
				r_v_buffer_e000_delay <= 0;
                r_v_buffer_000_delay <= 0;
                
				r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= 0;
				
				r_feedback_buffer <= 0;
				
                r_BRAM_read_buffer <= (r_cur_state == FWD_STBY)? r_BRAM_read_buffer:i_BRAM_read_data;
                r_waiting_buffer <= r_waiting_buffer;
				r_received_code_buffer <= r_received_code_buffer;
				o_c_message <= o_c_message;
			end
            FWD_FNLS: begin
			if (r_cur_state == FWD_FNLS) begin
				r_counter <= 0;
				
				r_v_buffer_e000_delay <= 0;
                r_v_buffer_000_delay <= 0;
                
				r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= 0;
				
				r_feedback_buffer <= 0;
				
                r_BRAM_read_buffer <= 0;
                r_waiting_buffer <= 0;
				r_received_code_buffer <= 0;
				o_c_message <= o_c_message;
				end
			else begin
				r_counter <= 0;
				
				r_v_buffer_e000_delay <= 0;
                r_v_buffer_000_delay <= 0;
                
				r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= 0;
				
				r_feedback_buffer <= 0;
				
                r_BRAM_read_buffer <= 0;
                r_waiting_buffer <= 0;
				r_received_code_buffer <= 0;
				o_c_message <= r_received_code_buffer;
				end
			end
			default: begin
				r_counter <= 0;
				
				r_v_buffer_e000_delay <= 0;
                r_v_buffer_000_delay <= 0;
                
				r_v_buffer_e000 <= 0;
				r_v_buffer_000 <= 0;
				
				r_feedback_buffer <= 0;
				
                r_BRAM_read_buffer <= 0;
                r_waiting_buffer <= 0;
				r_received_code_buffer <= 0;
				o_c_message <= 0;
			end
			endcase
	end
	
	
	
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// total: 8
	
	assign w_evaluated_term_S001_000[`D_CS_GF_ORDER -1:0] = w_ELP_term_000[`D_CS_GF_ORDER -1:0];
    assign w_evaluated_term_S002_000[`D_CS_GF_ORDER -1:0] = w_ELP_term_000[`D_CS_GF_ORDER -1:0];
    assign w_evaluated_term_S003_000[`D_CS_GF_ORDER -1:0] = w_ELP_term_000[`D_CS_GF_ORDER -1:0];
    assign w_evaluated_term_S004_000[`D_CS_GF_ORDER -1:0] = w_ELP_term_000[`D_CS_GF_ORDER -1:0];
    assign w_evaluated_term_S005_000[`D_CS_GF_ORDER -1:0] = w_ELP_term_000[`D_CS_GF_ORDER -1:0];
    assign w_evaluated_term_S006_000[`D_CS_GF_ORDER -1:0] = w_ELP_term_000[`D_CS_GF_ORDER -1:0];
    assign w_evaluated_term_S007_000[`D_CS_GF_ORDER -1:0] = w_ELP_term_000[`D_CS_GF_ORDER -1:0];
    assign w_evaluated_term_S008_000[`D_CS_GF_ORDER -1:0] = w_ELP_term_000[`D_CS_GF_ORDER -1:0];
	
	                                          ///
	                                        /////
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
	
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// total: 14

	d_CS_shortening_matrix_alpha_to_001 SM_001 ( // shortened by alpha_to_1879, 1879
    .i_in(r_v_buffer_e000[(  1+1)*`D_CS_GF_ORDER-1:(  1+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_001[`D_CS_GF_ORDER-1:0]) );

    d_CS_shortening_matrix_alpha_to_002 SM_002 ( // shortened by alpha_to_1879, 3758
    .i_in(r_v_buffer_e000[(  2+1)*`D_CS_GF_ORDER-1:(  2+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_002[`D_CS_GF_ORDER-1:0]) );

    d_CS_shortening_matrix_alpha_to_003 SM_003 ( // shortened by alpha_to_1879, 1542
    .i_in(r_v_buffer_e000[(  3+1)*`D_CS_GF_ORDER-1:(  3+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_003[`D_CS_GF_ORDER-1:0]) );

    d_CS_shortening_matrix_alpha_to_004 SM_004 ( // shortened by alpha_to_1879, 3421
    .i_in(r_v_buffer_e000[(  4+1)*`D_CS_GF_ORDER-1:(  4+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_004[`D_CS_GF_ORDER-1:0]) );

    d_CS_shortening_matrix_alpha_to_005 SM_005 ( // shortened by alpha_to_1879, 1205
    .i_in(r_v_buffer_e000[(  5+1)*`D_CS_GF_ORDER-1:(  5+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_005[`D_CS_GF_ORDER-1:0]) );

    d_CS_shortening_matrix_alpha_to_006 SM_006 ( // shortened by alpha_to_1879, 3084
    .i_in(r_v_buffer_e000[(  6+1)*`D_CS_GF_ORDER-1:(  6+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_006[`D_CS_GF_ORDER-1:0]) );

    d_CS_shortening_matrix_alpha_to_007 SM_007 ( // shortened by alpha_to_1879, 868
    .i_in(r_v_buffer_e000[(  7+1)*`D_CS_GF_ORDER-1:(  7+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_007[`D_CS_GF_ORDER-1:0]) );

    d_CS_shortening_matrix_alpha_to_008 SM_008 ( // shortened by alpha_to_1879, 2747
    .i_in(r_v_buffer_e000[(  8+1)*`D_CS_GF_ORDER-1:(  8+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_008[`D_CS_GF_ORDER-1:0]) );

    d_CS_shortening_matrix_alpha_to_009 SM_009 ( // shortened by alpha_to_1879, 531
    .i_in(r_v_buffer_e000[(  9+1)*`D_CS_GF_ORDER-1:(  9+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_009[`D_CS_GF_ORDER-1:0]) );

    d_CS_shortening_matrix_alpha_to_010 SM_010 ( // shortened by alpha_to_1879, 2410
    .i_in(r_v_buffer_e000[( 10+1)*`D_CS_GF_ORDER-1:( 10+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_010[`D_CS_GF_ORDER-1:0]) );

    d_CS_shortening_matrix_alpha_to_011 SM_011 ( // shortened by alpha_to_1879, 194
    .i_in(r_v_buffer_e000[( 11+1)*`D_CS_GF_ORDER-1:( 11+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_011[`D_CS_GF_ORDER-1:0]) );

    d_CS_shortening_matrix_alpha_to_012 SM_012 ( // shortened by alpha_to_1879, 2073
    .i_in(r_v_buffer_e000[( 12+1)*`D_CS_GF_ORDER-1:( 12+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_012[`D_CS_GF_ORDER-1:0]) );

    d_CS_shortening_matrix_alpha_to_013 SM_013 ( // shortened by alpha_to_1879, 3952
    .i_in(r_v_buffer_e000[( 13+1)*`D_CS_GF_ORDER-1:( 13+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_013[`D_CS_GF_ORDER-1:0]) );

    d_CS_shortening_matrix_alpha_to_014 SM_014 ( // shortened by alpha_to_1879, 1736
    .i_in(r_v_buffer_e000[( 14+1)*`D_CS_GF_ORDER-1:( 14+0)*`D_CS_GF_ORDER]), .o_out(w_shortened_v_014[`D_CS_GF_ORDER-1:0]) );
	                                         

											  ///
	                                        /////
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
	
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// total: 14 * 8 = 112
	
	d_CS_evaluation_matrix_slot_001_alpha_to_001 EM_S001_001 ( // evaluated by alpha_to_1, 1
    .i_in(w_ELP_term_001[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_001[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_001_alpha_to_002 EM_S001_002 ( // evaluated by alpha_to_1, 2
    .i_in(w_ELP_term_002[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_002[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_001_alpha_to_003 EM_S001_003 ( // evaluated by alpha_to_1, 3
    .i_in(w_ELP_term_003[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_003[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_001_alpha_to_004 EM_S001_004 ( // evaluated by alpha_to_1, 4
    .i_in(w_ELP_term_004[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_004[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_001_alpha_to_005 EM_S001_005 ( // evaluated by alpha_to_1, 5
    .i_in(w_ELP_term_005[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_005[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_001_alpha_to_006 EM_S001_006 ( // evaluated by alpha_to_1, 6
    .i_in(w_ELP_term_006[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_006[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_001_alpha_to_007 EM_S001_007 ( // evaluated by alpha_to_1, 7
    .i_in(w_ELP_term_007[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_007[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_001_alpha_to_008 EM_S001_008 ( // evaluated by alpha_to_1, 8
    .i_in(w_ELP_term_008[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_008[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_001_alpha_to_009 EM_S001_009 ( // evaluated by alpha_to_1, 9
    .i_in(w_ELP_term_009[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_009[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_001_alpha_to_010 EM_S001_010 ( // evaluated by alpha_to_1, 10
    .i_in(w_ELP_term_010[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_010[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_001_alpha_to_011 EM_S001_011 ( // evaluated by alpha_to_1, 11
    .i_in(w_ELP_term_011[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_011[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_001_alpha_to_012 EM_S001_012 ( // evaluated by alpha_to_1, 12
    .i_in(w_ELP_term_012[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_012[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_001_alpha_to_013 EM_S001_013 ( // evaluated by alpha_to_1, 13
    .i_in(w_ELP_term_013[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_013[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_001_alpha_to_014 EM_S001_014 ( // evaluated by alpha_to_1, 14
    .i_in(w_ELP_term_014[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S001_014[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_001 EM_S002_001 ( // evaluated by alpha_to_2, 2
    .i_in(w_ELP_term_001[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_001[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_002 EM_S002_002 ( // evaluated by alpha_to_2, 4
    .i_in(w_ELP_term_002[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_002[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_003 EM_S002_003 ( // evaluated by alpha_to_2, 6
    .i_in(w_ELP_term_003[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_003[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_004 EM_S002_004 ( // evaluated by alpha_to_2, 8
    .i_in(w_ELP_term_004[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_004[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_005 EM_S002_005 ( // evaluated by alpha_to_2, 10
    .i_in(w_ELP_term_005[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_005[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_006 EM_S002_006 ( // evaluated by alpha_to_2, 12
    .i_in(w_ELP_term_006[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_006[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_007 EM_S002_007 ( // evaluated by alpha_to_2, 14
    .i_in(w_ELP_term_007[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_007[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_008 EM_S002_008 ( // evaluated by alpha_to_2, 16
    .i_in(w_ELP_term_008[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_008[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_009 EM_S002_009 ( // evaluated by alpha_to_2, 18
    .i_in(w_ELP_term_009[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_009[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_010 EM_S002_010 ( // evaluated by alpha_to_2, 20
    .i_in(w_ELP_term_010[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_010[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_011 EM_S002_011 ( // evaluated by alpha_to_2, 22
    .i_in(w_ELP_term_011[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_011[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_012 EM_S002_012 ( // evaluated by alpha_to_2, 24
    .i_in(w_ELP_term_012[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_012[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_013 EM_S002_013 ( // evaluated by alpha_to_2, 26
    .i_in(w_ELP_term_013[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_013[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_002_alpha_to_014 EM_S002_014 ( // evaluated by alpha_to_2, 28
    .i_in(w_ELP_term_014[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S002_014[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_001 EM_S003_001 ( // evaluated by alpha_to_3, 3
    .i_in(w_ELP_term_001[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_001[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_002 EM_S003_002 ( // evaluated by alpha_to_3, 6
    .i_in(w_ELP_term_002[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_002[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_003 EM_S003_003 ( // evaluated by alpha_to_3, 9
    .i_in(w_ELP_term_003[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_003[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_004 EM_S003_004 ( // evaluated by alpha_to_3, 12
    .i_in(w_ELP_term_004[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_004[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_005 EM_S003_005 ( // evaluated by alpha_to_3, 15
    .i_in(w_ELP_term_005[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_005[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_006 EM_S003_006 ( // evaluated by alpha_to_3, 18
    .i_in(w_ELP_term_006[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_006[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_007 EM_S003_007 ( // evaluated by alpha_to_3, 21
    .i_in(w_ELP_term_007[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_007[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_008 EM_S003_008 ( // evaluated by alpha_to_3, 24
    .i_in(w_ELP_term_008[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_008[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_009 EM_S003_009 ( // evaluated by alpha_to_3, 27
    .i_in(w_ELP_term_009[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_009[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_010 EM_S003_010 ( // evaluated by alpha_to_3, 30
    .i_in(w_ELP_term_010[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_010[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_011 EM_S003_011 ( // evaluated by alpha_to_3, 33
    .i_in(w_ELP_term_011[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_011[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_012 EM_S003_012 ( // evaluated by alpha_to_3, 36
    .i_in(w_ELP_term_012[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_012[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_013 EM_S003_013 ( // evaluated by alpha_to_3, 39
    .i_in(w_ELP_term_013[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_013[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_003_alpha_to_014 EM_S003_014 ( // evaluated by alpha_to_3, 42
    .i_in(w_ELP_term_014[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S003_014[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_001 EM_S004_001 ( // evaluated by alpha_to_4, 4
    .i_in(w_ELP_term_001[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_001[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_002 EM_S004_002 ( // evaluated by alpha_to_4, 8
    .i_in(w_ELP_term_002[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_002[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_003 EM_S004_003 ( // evaluated by alpha_to_4, 12
    .i_in(w_ELP_term_003[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_003[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_004 EM_S004_004 ( // evaluated by alpha_to_4, 16
    .i_in(w_ELP_term_004[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_004[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_005 EM_S004_005 ( // evaluated by alpha_to_4, 20
    .i_in(w_ELP_term_005[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_005[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_006 EM_S004_006 ( // evaluated by alpha_to_4, 24
    .i_in(w_ELP_term_006[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_006[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_007 EM_S004_007 ( // evaluated by alpha_to_4, 28
    .i_in(w_ELP_term_007[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_007[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_008 EM_S004_008 ( // evaluated by alpha_to_4, 32
    .i_in(w_ELP_term_008[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_008[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_009 EM_S004_009 ( // evaluated by alpha_to_4, 36
    .i_in(w_ELP_term_009[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_009[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_010 EM_S004_010 ( // evaluated by alpha_to_4, 40
    .i_in(w_ELP_term_010[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_010[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_011 EM_S004_011 ( // evaluated by alpha_to_4, 44
    .i_in(w_ELP_term_011[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_011[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_012 EM_S004_012 ( // evaluated by alpha_to_4, 48
    .i_in(w_ELP_term_012[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_012[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_013 EM_S004_013 ( // evaluated by alpha_to_4, 52
    .i_in(w_ELP_term_013[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_013[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_004_alpha_to_014 EM_S004_014 ( // evaluated by alpha_to_4, 56
    .i_in(w_ELP_term_014[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S004_014[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_001 EM_S005_001 ( // evaluated by alpha_to_5, 5
    .i_in(w_ELP_term_001[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_001[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_002 EM_S005_002 ( // evaluated by alpha_to_5, 10
    .i_in(w_ELP_term_002[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_002[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_003 EM_S005_003 ( // evaluated by alpha_to_5, 15
    .i_in(w_ELP_term_003[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_003[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_004 EM_S005_004 ( // evaluated by alpha_to_5, 20
    .i_in(w_ELP_term_004[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_004[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_005 EM_S005_005 ( // evaluated by alpha_to_5, 25
    .i_in(w_ELP_term_005[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_005[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_006 EM_S005_006 ( // evaluated by alpha_to_5, 30
    .i_in(w_ELP_term_006[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_006[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_007 EM_S005_007 ( // evaluated by alpha_to_5, 35
    .i_in(w_ELP_term_007[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_007[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_008 EM_S005_008 ( // evaluated by alpha_to_5, 40
    .i_in(w_ELP_term_008[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_008[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_009 EM_S005_009 ( // evaluated by alpha_to_5, 45
    .i_in(w_ELP_term_009[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_009[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_010 EM_S005_010 ( // evaluated by alpha_to_5, 50
    .i_in(w_ELP_term_010[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_010[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_011 EM_S005_011 ( // evaluated by alpha_to_5, 55
    .i_in(w_ELP_term_011[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_011[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_012 EM_S005_012 ( // evaluated by alpha_to_5, 60
    .i_in(w_ELP_term_012[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_012[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_013 EM_S005_013 ( // evaluated by alpha_to_5, 65
    .i_in(w_ELP_term_013[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_013[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_005_alpha_to_014 EM_S005_014 ( // evaluated by alpha_to_5, 70
    .i_in(w_ELP_term_014[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S005_014[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_001 EM_S006_001 ( // evaluated by alpha_to_6, 6
    .i_in(w_ELP_term_001[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_001[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_002 EM_S006_002 ( // evaluated by alpha_to_6, 12
    .i_in(w_ELP_term_002[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_002[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_003 EM_S006_003 ( // evaluated by alpha_to_6, 18
    .i_in(w_ELP_term_003[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_003[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_004 EM_S006_004 ( // evaluated by alpha_to_6, 24
    .i_in(w_ELP_term_004[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_004[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_005 EM_S006_005 ( // evaluated by alpha_to_6, 30
    .i_in(w_ELP_term_005[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_005[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_006 EM_S006_006 ( // evaluated by alpha_to_6, 36
    .i_in(w_ELP_term_006[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_006[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_007 EM_S006_007 ( // evaluated by alpha_to_6, 42
    .i_in(w_ELP_term_007[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_007[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_008 EM_S006_008 ( // evaluated by alpha_to_6, 48
    .i_in(w_ELP_term_008[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_008[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_009 EM_S006_009 ( // evaluated by alpha_to_6, 54
    .i_in(w_ELP_term_009[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_009[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_010 EM_S006_010 ( // evaluated by alpha_to_6, 60
    .i_in(w_ELP_term_010[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_010[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_011 EM_S006_011 ( // evaluated by alpha_to_6, 66
    .i_in(w_ELP_term_011[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_011[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_012 EM_S006_012 ( // evaluated by alpha_to_6, 72
    .i_in(w_ELP_term_012[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_012[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_013 EM_S006_013 ( // evaluated by alpha_to_6, 78
    .i_in(w_ELP_term_013[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_013[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_006_alpha_to_014 EM_S006_014 ( // evaluated by alpha_to_6, 84
    .i_in(w_ELP_term_014[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S006_014[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_001 EM_S007_001 ( // evaluated by alpha_to_7, 7
    .i_in(w_ELP_term_001[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_001[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_002 EM_S007_002 ( // evaluated by alpha_to_7, 14
    .i_in(w_ELP_term_002[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_002[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_003 EM_S007_003 ( // evaluated by alpha_to_7, 21
    .i_in(w_ELP_term_003[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_003[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_004 EM_S007_004 ( // evaluated by alpha_to_7, 28
    .i_in(w_ELP_term_004[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_004[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_005 EM_S007_005 ( // evaluated by alpha_to_7, 35
    .i_in(w_ELP_term_005[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_005[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_006 EM_S007_006 ( // evaluated by alpha_to_7, 42
    .i_in(w_ELP_term_006[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_006[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_007 EM_S007_007 ( // evaluated by alpha_to_7, 49
    .i_in(w_ELP_term_007[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_007[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_008 EM_S007_008 ( // evaluated by alpha_to_7, 56
    .i_in(w_ELP_term_008[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_008[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_009 EM_S007_009 ( // evaluated by alpha_to_7, 63
    .i_in(w_ELP_term_009[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_009[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_010 EM_S007_010 ( // evaluated by alpha_to_7, 70
    .i_in(w_ELP_term_010[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_010[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_011 EM_S007_011 ( // evaluated by alpha_to_7, 77
    .i_in(w_ELP_term_011[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_011[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_012 EM_S007_012 ( // evaluated by alpha_to_7, 84
    .i_in(w_ELP_term_012[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_012[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_013 EM_S007_013 ( // evaluated by alpha_to_7, 91
    .i_in(w_ELP_term_013[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_013[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_007_alpha_to_014 EM_S007_014 ( // evaluated by alpha_to_7, 98
    .i_in(w_ELP_term_014[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S007_014[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_001 EM_S008_001 ( // evaluated by alpha_to_8, 8
    .i_in(w_ELP_term_001[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_001[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_002 EM_S008_002 ( // evaluated by alpha_to_8, 16
    .i_in(w_ELP_term_002[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_002[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_003 EM_S008_003 ( // evaluated by alpha_to_8, 24
    .i_in(w_ELP_term_003[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_003[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_004 EM_S008_004 ( // evaluated by alpha_to_8, 32
    .i_in(w_ELP_term_004[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_004[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_005 EM_S008_005 ( // evaluated by alpha_to_8, 40
    .i_in(w_ELP_term_005[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_005[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_006 EM_S008_006 ( // evaluated by alpha_to_8, 48
    .i_in(w_ELP_term_006[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_006[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_007 EM_S008_007 ( // evaluated by alpha_to_8, 56
    .i_in(w_ELP_term_007[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_007[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_008 EM_S008_008 ( // evaluated by alpha_to_8, 64
    .i_in(w_ELP_term_008[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_008[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_009 EM_S008_009 ( // evaluated by alpha_to_8, 72
    .i_in(w_ELP_term_009[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_009[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_010 EM_S008_010 ( // evaluated by alpha_to_8, 80
    .i_in(w_ELP_term_010[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_010[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_011 EM_S008_011 ( // evaluated by alpha_to_8, 88
    .i_in(w_ELP_term_011[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_011[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_012 EM_S008_012 ( // evaluated by alpha_to_8, 96
    .i_in(w_ELP_term_012[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_012[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_013 EM_S008_013 ( // evaluated by alpha_to_8, 104
    .i_in(w_ELP_term_013[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_013[`D_CS_GF_ORDER-1:0]) );

    d_CS_evaluation_matrix_slot_008_alpha_to_014 EM_S008_014 ( // evaluated by alpha_to_8, 112
    .i_in(w_ELP_term_014[`D_CS_GF_ORDER-1:0]), .o_out(w_evaluated_term_S008_014[`D_CS_GF_ORDER-1:0]) );
	
	                                          ///
	                                        /////
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
	
	/////////////////////////////////////////////
	////////// GENERATED BY C PROGRAMA //////////
	/////
	///
	
	// total: 8, 8, 1
	
	assign w_slot_001_flip = |( w_evaluated_term_S001_000[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_001[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_002[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_003[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_004[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_005[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_006[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_007[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_008[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_009[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_010[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_011[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_012[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_013[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S001_014[`D_CS_GF_ORDER-1:0] );
    assign w_slot_002_flip = |( w_evaluated_term_S002_000[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_001[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_002[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_003[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_004[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_005[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_006[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_007[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_008[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_009[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_010[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_011[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_012[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_013[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S002_014[`D_CS_GF_ORDER-1:0] );
    assign w_slot_003_flip = |( w_evaluated_term_S003_000[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_001[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_002[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_003[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_004[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_005[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_006[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_007[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_008[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_009[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_010[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_011[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_012[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_013[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S003_014[`D_CS_GF_ORDER-1:0] );
    assign w_slot_004_flip = |( w_evaluated_term_S004_000[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_001[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_002[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_003[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_004[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_005[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_006[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_007[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_008[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_009[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_010[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_011[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_012[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_013[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S004_014[`D_CS_GF_ORDER-1:0] );
    assign w_slot_005_flip = |( w_evaluated_term_S005_000[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_001[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_002[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_003[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_004[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_005[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_006[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_007[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_008[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_009[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_010[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_011[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_012[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_013[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S005_014[`D_CS_GF_ORDER-1:0] );
    assign w_slot_006_flip = |( w_evaluated_term_S006_000[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_001[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_002[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_003[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_004[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_005[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_006[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_007[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_008[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_009[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_010[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_011[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_012[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_013[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S006_014[`D_CS_GF_ORDER-1:0] );
    assign w_slot_007_flip = |( w_evaluated_term_S007_000[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_001[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_002[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_003[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_004[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_005[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_006[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_007[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_008[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_009[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_010[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_011[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_012[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_013[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S007_014[`D_CS_GF_ORDER-1:0] );
    assign w_slot_008_flip = |( w_evaluated_term_S008_000[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_001[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_002[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_003[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_004[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_005[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_006[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_007[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_008[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_009[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_010[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_011[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_012[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_013[`D_CS_GF_ORDER-1:0] ^ w_evaluated_term_S008_014[`D_CS_GF_ORDER-1:0] );

    assign w_slot_001_flipped_message = ~( w_slot_001_flip ^ r_received_code_buffer[7] );
    assign w_slot_002_flipped_message = ~( w_slot_002_flip ^ r_received_code_buffer[6] );
    assign w_slot_003_flipped_message = ~( w_slot_003_flip ^ r_received_code_buffer[5] );
    assign w_slot_004_flipped_message = ~( w_slot_004_flip ^ r_received_code_buffer[4] );
    assign w_slot_005_flipped_message = ~( w_slot_005_flip ^ r_received_code_buffer[3] );
    assign w_slot_006_flipped_message = ~( w_slot_006_flip ^ r_received_code_buffer[2] );
    assign w_slot_007_flipped_message = ~( w_slot_007_flip ^ r_received_code_buffer[1] );
    assign w_slot_008_flipped_message = ~( w_slot_008_flip ^ r_received_code_buffer[0] );

    assign w_flipped_message[`D_CS_P_LVL-1:0] = { w_slot_001_flipped_message, w_slot_002_flipped_message, w_slot_003_flipped_message, w_slot_004_flipped_message, w_slot_005_flipped_message, w_slot_006_flipped_message, w_slot_007_flipped_message, w_slot_008_flipped_message };
	
	                                          ///
	                                        /////
	////////// GENERATED BY C PROGRAMA //////////
	/////////////////////////////////////////////
	
endmodule
