

`timescale 1ns / 1ps

module SCFIFO_40x64_withCount
(
    input           iClock          ,
    input           iReset          ,

    input   [39:0]  iPushData       ,
    input           iPushEnable     ,
    output          oIsFull         ,
    
    output  [39:0]  oPopData        ,
    input           iPopEnable      ,
    output          oIsEmpty        ,
    
    output  [5:0]   oDataCount
);

  wire [6:0] data_count_internal;

    SCFIFO_sync #(
        .DATA_WIDTH(40),
        .FIFO_DEPTH(64)
    ) u1_fifo_sync (
        .clk        (iClock),
        .rst        (iReset),
        .wr_en      (iPushEnable),
        .wr_data    (iPushData),
        .wr_full    (oIsFull),
        .rd_en      (iPopEnable),
        .rd_data    (oPopData),
        .rd_empty   (oIsEmpty),
        .data_count (data_count_internal)
    );
assign oDataCount = data_count_internal[5:0];


endmodule
