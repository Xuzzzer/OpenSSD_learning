


`define D_CS_GF_ORDER 12 // Galois field order, GF(2^12)
`define D_CS_ECC_T 14 // error correction capability t = 14

`define D_CS_P_LVL 8 // data area BCH decoder CS parallel level

`define D_CS_O_CNT 256 // no corrected parity output, 256B chunk / 8b = 256
`define D_CS_O_CNT_BIT 9 // bigger than CS_OUTPUT_LOOP_COUNT, 2^8 = 256
