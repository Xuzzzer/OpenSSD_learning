

`timescale 1ns / 1ps


module dma_if # (
	parameter 	P_SLOT_TAG_WIDTH			=  10, //slot_modified
	parameter	C_PCIE_DATA_WIDTH			= 512,
	parameter	C_PCIE_ADDR_WIDTH			= 48, //modified
	parameter	C_M_AXI_DATA_WIDTH			= 64
)
(
	input									pcie_user_clk,
	input									pcie_user_rst_n,

	input	[1:0]							pcie_max_payload_size,
	input	[2:0]							pcie_max_read_req_size,
	input									pcie_rcb,

	output	[(P_SLOT_TAG_WIDTH+1)-1:0]		hcmd_prp_rd_addr,//slot_modified
	input	[53:0]							hcmd_prp_rd_data, //modified

	output									hcmd_nlb_wr1_en, 
	output	[P_SLOT_TAG_WIDTH-1:0]			hcmd_nlb_wr1_addr,//slot_modified
	output	[18:0]							hcmd_nlb_wr1_data,
	input									hcmd_nlb_wr1_rdy_n,

	output	[P_SLOT_TAG_WIDTH-1:0]			hcmd_nlb_rd_addr, //slot_modified
	input	[18:0]							hcmd_nlb_rd_data,

	output									dev_rx_cmd_wr_en,
	output	[29:0]							dev_rx_cmd_wr_data,
	input									dev_rx_cmd_full_n,

	output									dev_tx_cmd_wr_en,
	output	[29:0]							dev_tx_cmd_wr_data,
	input									dev_tx_cmd_full_n,

	output									tx_prp_mrd_req,
	output	[7:0]							tx_prp_mrd_tag,
	output	[12:2]							tx_prp_mrd_len,
	output	[C_PCIE_ADDR_WIDTH-1:2]			tx_prp_mrd_addr,
	input									tx_prp_mrd_req_ack,

	input	[7:0]							cpld_prp_fifo_tag,
	input	[C_PCIE_DATA_WIDTH-1:0]			cpld_prp_fifo_wr_data,
	input									cpld_prp_fifo_wr_en,
	input									cpld_prp_fifo_tag_last,

	output									tx_dma_mrd_req,
	output	[7:0]							tx_dma_mrd_tag,
	output	[12:2]							tx_dma_mrd_len,
	output	[C_PCIE_ADDR_WIDTH-1:2]			tx_dma_mrd_addr,
	input									tx_dma_mrd_req_ack,

	input	[7:0]							cpld_dma_fifo_tag,
	input	[C_PCIE_DATA_WIDTH-1:0]			cpld_dma_fifo_wr_data,
	input									cpld_dma_fifo_wr_en,
	input									cpld_dma_fifo_tag_last,

	output									tx_dma_mwr_req,
	output	[7:0]							tx_dma_mwr_tag,
	output	[12:2]							tx_dma_mwr_len,
	output	[C_PCIE_ADDR_WIDTH-1:2]			tx_dma_mwr_addr,
	input									tx_dma_mwr_req_ack,
	input									tx_dma_mwr_data_last,

	input									pcie_tx_dma_fifo_rd_en,
	output	[C_PCIE_DATA_WIDTH-1:0]			pcie_tx_dma_fifo_rd_data,

	output									hcmd_cq_wr0_en,
	output	[(P_SLOT_TAG_WIDTH+28)-1:0]		hcmd_cq_wr0_data0, //slot_modified
	output	[(P_SLOT_TAG_WIDTH+28)-1:0]		hcmd_cq_wr0_data1, //slot_modified
	input									hcmd_cq_wr0_rdy_n,

	input									cpu_bus_clk,
	input									cpu_bus_rst_n,

	input									dma_cmd_wr_en,
	input	[55:0]							dma_cmd_wr_data0, //modified
	input	[55:0]							dma_cmd_wr_data1, //modified
	output									dma_cmd_wr_rdy_n,

	output	[7:0]							dma_rx_direct_done_cnt,
	output	[7:0]							dma_tx_direct_done_cnt,
	output	[7:0]							dma_rx_done_cnt,
	output	[7:0]							dma_tx_done_cnt,

	input									dma_bus_clk,
	input									dma_bus_rst_n,

	input									pcie_rx_fifo_rd_en,
	output	[C_M_AXI_DATA_WIDTH-1:0]		pcie_rx_fifo_rd_data,
	input									pcie_rx_fifo_free_en,
	input	[10:6]							pcie_rx_fifo_free_len, 
	output									pcie_rx_fifo_empty_n,

	input									pcie_tx_fifo_alloc_en,
	input	[10:6]							pcie_tx_fifo_alloc_len, 
	input									pcie_tx_fifo_wr_en,
	input	[C_M_AXI_DATA_WIDTH-1:0]		pcie_tx_fifo_wr_data,
	output									pcie_tx_fifo_full_n,

	input									dma_rx_done_wr_en,
	input	[(P_SLOT_TAG_WIDTH+15)-1:0]		dma_rx_done_wr_data, //slot_modified
	output									dma_rx_done_wr_rdy_n
);

wire										w_pcie_rx_cmd_wr_en;
wire	[45:0]								w_pcie_rx_cmd_wr_data; //modified
wire										w_pcie_rx_cmd_full_n;

wire										w_pcie_tx_cmd_wr_en;
wire	[45:0]								w_pcie_tx_cmd_wr_data; //modified
wire										w_pcie_tx_cmd_full_n;

wire										w_dma_tx_done_wr_en;
wire	[(P_SLOT_TAG_WIDTH+15)-1:0]			w_dma_tx_done_wr_data; //slot_modified
wire										w_dma_tx_done_wr_rdy_n;


dma_cmd # (
	.P_SLOT_TAG_WIDTH						(P_SLOT_TAG_WIDTH) //slot_modified
)
dma_cmd_inst0
(
	.pcie_user_clk							(pcie_user_clk),
	.pcie_user_rst_n						(pcie_user_rst_n),

	.pcie_rcb								(pcie_rcb),

	.hcmd_prp_rd_addr						(hcmd_prp_rd_addr),
	.hcmd_prp_rd_data						(hcmd_prp_rd_data),

	.hcmd_nlb_wr1_en						(hcmd_nlb_wr1_en),
	.hcmd_nlb_wr1_addr						(hcmd_nlb_wr1_addr),
	.hcmd_nlb_wr1_data						(hcmd_nlb_wr1_data),
	.hcmd_nlb_wr1_rdy_n						(hcmd_nlb_wr1_rdy_n),

	.hcmd_nlb_rd_addr						(hcmd_nlb_rd_addr),
	.hcmd_nlb_rd_data						(hcmd_nlb_rd_data),

	.dev_rx_cmd_wr_en						(dev_rx_cmd_wr_en),
	.dev_rx_cmd_wr_data						(dev_rx_cmd_wr_data),
	.dev_rx_cmd_full_n						(dev_rx_cmd_full_n),

	.dev_tx_cmd_wr_en						(dev_tx_cmd_wr_en),
	.dev_tx_cmd_wr_data						(dev_tx_cmd_wr_data),
	.dev_tx_cmd_full_n						(dev_tx_cmd_full_n),

	.tx_prp_mrd_req							(tx_prp_mrd_req),
	.tx_prp_mrd_tag							(tx_prp_mrd_tag),
	.tx_prp_mrd_len							(tx_prp_mrd_len),
	.tx_prp_mrd_addr						(tx_prp_mrd_addr),
	.tx_prp_mrd_req_ack						(tx_prp_mrd_req_ack),

	.cpld_prp_fifo_tag						(cpld_prp_fifo_tag),
	.cpld_prp_fifo_wr_data					(cpld_prp_fifo_wr_data),
	.cpld_prp_fifo_wr_en					(cpld_prp_fifo_wr_en),
	.cpld_prp_fifo_tag_last					(cpld_prp_fifo_tag_last),

	.pcie_rx_cmd_wr_en						(w_pcie_rx_cmd_wr_en),
	.pcie_rx_cmd_wr_data					(w_pcie_rx_cmd_wr_data),
	.pcie_rx_cmd_full_n						(w_pcie_rx_cmd_full_n),

	.pcie_tx_cmd_wr_en						(w_pcie_tx_cmd_wr_en),
	.pcie_tx_cmd_wr_data					(w_pcie_tx_cmd_wr_data),
	.pcie_tx_cmd_full_n						(w_pcie_tx_cmd_full_n),

	.dma_tx_done_wr_en						(w_dma_tx_done_wr_en),
	.dma_tx_done_wr_data					(w_dma_tx_done_wr_data),
	.dma_tx_done_wr_rdy_n					(w_dma_tx_done_wr_rdy_n),

	.hcmd_cq_wr0_en							(hcmd_cq_wr0_en),
	.hcmd_cq_wr0_data0						(hcmd_cq_wr0_data0),
	.hcmd_cq_wr0_data1						(hcmd_cq_wr0_data1),
	.hcmd_cq_wr0_rdy_n						(hcmd_cq_wr0_rdy_n),

	.cpu_bus_clk							(cpu_bus_clk),
	.cpu_bus_rst_n							(cpu_bus_rst_n),

	.dma_cmd_wr_en							(dma_cmd_wr_en),
	.dma_cmd_wr_data0						(dma_cmd_wr_data0),
	.dma_cmd_wr_data1						(dma_cmd_wr_data1),
	.dma_cmd_wr_rdy_n						(dma_cmd_wr_rdy_n),

	.dma_rx_direct_done_cnt					(dma_rx_direct_done_cnt),
	.dma_tx_direct_done_cnt					(dma_tx_direct_done_cnt),
	.dma_rx_done_cnt						(dma_rx_done_cnt),
	.dma_tx_done_cnt						(dma_tx_done_cnt),

	.dma_bus_clk							(dma_bus_clk),
	.dma_bus_rst_n							(dma_bus_rst_n),

	.dma_rx_done_wr_en						(dma_rx_done_wr_en),
	.dma_rx_done_wr_data					(dma_rx_done_wr_data),
	.dma_rx_done_wr_rdy_n					(dma_rx_done_wr_rdy_n)
);

pcie_rx_dma
pcie_rx_dma_inst0
(
	.pcie_user_clk							(pcie_user_clk),
	.pcie_user_rst_n						(pcie_user_rst_n),

	.pcie_max_read_req_size					(pcie_max_read_req_size),

	.pcie_rx_cmd_wr_en						(w_pcie_rx_cmd_wr_en),
	.pcie_rx_cmd_wr_data					(w_pcie_rx_cmd_wr_data),
	.pcie_rx_cmd_full_n						(w_pcie_rx_cmd_full_n),

	.tx_dma_mrd_req							(tx_dma_mrd_req),
	.tx_dma_mrd_tag							(tx_dma_mrd_tag),
	.tx_dma_mrd_len							(tx_dma_mrd_len),
	.tx_dma_mrd_addr						(tx_dma_mrd_addr),
	.tx_dma_mrd_req_ack						(tx_dma_mrd_req_ack),

	.cpld_dma_fifo_tag						(cpld_dma_fifo_tag),
	.cpld_dma_fifo_wr_data					(cpld_dma_fifo_wr_data),
	.cpld_dma_fifo_wr_en					(cpld_dma_fifo_wr_en),
	.cpld_dma_fifo_tag_last					(cpld_dma_fifo_tag_last),

	.dma_bus_clk							(dma_bus_clk),
	.dma_bus_rst_n							(dma_bus_rst_n),

	.pcie_rx_fifo_rd_en						(pcie_rx_fifo_rd_en),
	.pcie_rx_fifo_rd_data					(pcie_rx_fifo_rd_data),
	.pcie_rx_fifo_free_en					(pcie_rx_fifo_free_en),
	.pcie_rx_fifo_free_len					(pcie_rx_fifo_free_len),
	.pcie_rx_fifo_empty_n					(pcie_rx_fifo_empty_n)
);

pcie_tx_dma # (
	.P_SLOT_TAG_WIDTH						(P_SLOT_TAG_WIDTH) //slot_modified
)
pcie_tx_dma_inst0
(
	.pcie_user_clk							(pcie_user_clk),
	.pcie_user_rst_n						(pcie_user_rst_n),

	.pcie_max_payload_size					(pcie_max_payload_size),

	.pcie_tx_cmd_wr_en						(w_pcie_tx_cmd_wr_en),
	.pcie_tx_cmd_wr_data					(w_pcie_tx_cmd_wr_data),
	.pcie_tx_cmd_full_n						(w_pcie_tx_cmd_full_n),

	.tx_dma_mwr_req							(tx_dma_mwr_req),
	.tx_dma_mwr_tag							(tx_dma_mwr_tag),
	.tx_dma_mwr_len							(tx_dma_mwr_len),
	.tx_dma_mwr_addr						(tx_dma_mwr_addr),
	.tx_dma_mwr_req_ack						(tx_dma_mwr_req_ack),
	.tx_dma_mwr_data_last					(tx_dma_mwr_data_last),

	.pcie_tx_dma_fifo_rd_en					(pcie_tx_dma_fifo_rd_en),
	.pcie_tx_dma_fifo_rd_data				(pcie_tx_dma_fifo_rd_data),

	.dma_tx_done_wr_en						(w_dma_tx_done_wr_en),
	.dma_tx_done_wr_data					(w_dma_tx_done_wr_data),
	.dma_tx_done_wr_rdy_n					(w_dma_tx_done_wr_rdy_n),

	.dma_bus_clk							(dma_bus_clk),
	.dma_bus_rst_n							(dma_bus_rst_n),

	.pcie_tx_fifo_alloc_en					(pcie_tx_fifo_alloc_en),
	.pcie_tx_fifo_alloc_len					(pcie_tx_fifo_alloc_len),
	.pcie_tx_fifo_wr_en						(pcie_tx_fifo_wr_en),
	.pcie_tx_fifo_wr_data					(pcie_tx_fifo_wr_data),
	.pcie_tx_fifo_full_n					(pcie_tx_fifo_full_n)
);

endmodule
