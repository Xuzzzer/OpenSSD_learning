


`timescale 1ns / 1ps

module pcie_hcmd # (
	parameter	C_PCIE_DATA_WIDTH			= 512,
	parameter	C_PCIE_ADDR_WIDTH			= 48, //modified
	parameter 	P_SLOT_TAG_WIDTH			=  10, //slot_modified
	parameter 	P_SLOT_WIDTH				= 1024 //slot_modified
)
(
	input									pcie_user_clk,
	input									pcie_user_rst_n,

	input	[C_PCIE_ADDR_WIDTH-1:2]			admin_sq_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			admin_cq_bs_addr,
	input	[7:0]							admin_sq_size,
	input	[7:0]							admin_cq_size,

	input	[7:0]							admin_sq_tail_ptr,
	input	[7:0]							io_sq1_tail_ptr,
	input	[7:0]							io_sq2_tail_ptr,
	input	[7:0]							io_sq3_tail_ptr,
	input	[7:0]							io_sq4_tail_ptr,
	input	[7:0]							io_sq5_tail_ptr,
	input	[7:0]							io_sq6_tail_ptr,
	input	[7:0]							io_sq7_tail_ptr,
	input	[7:0]							io_sq8_tail_ptr,

	input	[7:0]							cpld_sq_fifo_tag,
	input	[C_PCIE_DATA_WIDTH-1:0]			cpld_sq_fifo_wr_data,
	input									cpld_sq_fifo_wr_en,
	input									cpld_sq_fifo_tag_last,

	output									tx_mrd_req,
	output	[7:0]							tx_mrd_tag,
	output	[12:2]							tx_mrd_len,
	output	[C_PCIE_ADDR_WIDTH-1:2]			tx_mrd_addr,
	input									tx_mrd_req_ack,

	output	[7:0]							admin_cq_tail_ptr,
	output	[7:0]							io_cq1_tail_ptr,
	output	[7:0]							io_cq2_tail_ptr,
	output	[7:0]							io_cq3_tail_ptr,
	output	[7:0]							io_cq4_tail_ptr,
	output	[7:0]							io_cq5_tail_ptr,
	output	[7:0]							io_cq6_tail_ptr,
	output	[7:0]							io_cq7_tail_ptr,
	output	[7:0]							io_cq8_tail_ptr,

	output									tx_cq_mwr_req,
	output	[7:0]							tx_cq_mwr_tag,
	output	[12:2]							tx_cq_mwr_len,
	output	[C_PCIE_ADDR_WIDTH-1:2]			tx_cq_mwr_addr,
	input									tx_cq_mwr_req_ack,
	input									tx_cq_mwr_rd_en,
	output	[C_PCIE_DATA_WIDTH-1:0]			tx_cq_mwr_rd_data,
	input									tx_cq_mwr_data_last,

	input	[(P_SLOT_TAG_WIDTH+1)-1:0]		hcmd_prp_rd_addr, //slot_modified
	output	[53:0]							hcmd_prp_rd_data, //modified

	input									hcmd_nlb_wr1_en,
	input	[P_SLOT_TAG_WIDTH-1:0]			hcmd_nlb_wr1_addr, //slot_modified
	input	[18:0]							hcmd_nlb_wr1_data,
	output									hcmd_nlb_wr1_rdy_n,

	input	[P_SLOT_TAG_WIDTH-1:0]			hcmd_nlb_rd_addr, //slot_modified
	output	[18:0]							hcmd_nlb_rd_data,

	input									hcmd_cq_wr0_en,
	input	[(P_SLOT_TAG_WIDTH+28)-1:0]		hcmd_cq_wr0_data0, //slot_modified
	input	[(P_SLOT_TAG_WIDTH+28)-1:0]		hcmd_cq_wr0_data1, //slot_modified
	output									hcmd_cq_wr0_rdy_n,
	
	input									cpu_bus_clk,
	input									cpu_bus_rst_n,

	input	[8:0]							sq_rst_n,
	input	[8:0]							sq_valid,
	input	[7:0]							io_sq1_size,
	input	[7:0]							io_sq2_size,
	input	[7:0]							io_sq3_size,
	input	[7:0]							io_sq4_size,
	input	[7:0]							io_sq5_size,
	input	[7:0]							io_sq6_size,
	input	[7:0]							io_sq7_size,
	input	[7:0]							io_sq8_size,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq1_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq2_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq3_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq4_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq5_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq6_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq7_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq8_bs_addr,
	input	[3:0]							io_sq1_cq_vec,
	input	[3:0]							io_sq2_cq_vec,
	input	[3:0]							io_sq3_cq_vec,
	input	[3:0]							io_sq4_cq_vec,
	input	[3:0]							io_sq5_cq_vec,
	input	[3:0]							io_sq6_cq_vec,
	input	[3:0]							io_sq7_cq_vec,
	input	[3:0]							io_sq8_cq_vec,

	input	[8:0]							cq_rst_n,
	input	[8:0]							cq_valid,
	input	[7:0]							io_cq1_size,
	input	[7:0]							io_cq2_size,
	input	[7:0]							io_cq3_size,
	input	[7:0]							io_cq4_size,
	input	[7:0]							io_cq5_size,
	input	[7:0]							io_cq6_size,
	input	[7:0]							io_cq7_size,
	input	[7:0]							io_cq8_size,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_cq1_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_cq2_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_cq3_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_cq4_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_cq5_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_cq6_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_cq7_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_cq8_bs_addr,

	input									hcmd_sq_rd_en,
	output	[(P_SLOT_TAG_WIDTH+12)-1:0]		hcmd_sq_rd_data,  //slot_modified
	output									hcmd_sq_empty_n,

	input	[(P_SLOT_TAG_WIDTH+2)+1:0]		hcmd_table_rd_addr, //slot_modified
	output	[31:0]							hcmd_table_rd_data,

	input									hcmd_cq_wr1_en,
	input	[(P_SLOT_TAG_WIDTH+28)-1:0]		hcmd_cq_wr1_data0,//slot_modified
	input	[(P_SLOT_TAG_WIDTH+28)-1:0]		hcmd_cq_wr1_data1,//slot_modified
	output									hcmd_cq_wr1_rdy_n
);

wire										w_hcmd_table_wr_en;
wire	[(P_SLOT_TAG_WIDTH+2)-1:0]			w_hcmd_table_wr_addr; //slot_modified
wire	[127:0]								w_hcmd_table_wr_data;

wire										w_hcmd_cid_wr_en;
wire	[P_SLOT_TAG_WIDTH-1:0]				w_hcmd_cid_wr_addr; //slot_modified
wire	[19:0]								w_hcmd_cid_wr_data;

wire	[P_SLOT_TAG_WIDTH-1:0]				w_hcmd_cid_rd_addr; //slot_modified
wire	[19:0]								w_hcmd_cid_rd_data;

wire										w_hcmd_prp_wr_en;
wire	[(P_SLOT_TAG_WIDTH+1)-1:0]			w_hcmd_prp_wr_addr; //slot_modified
wire	[53:0]								w_hcmd_prp_wr_data; //modified

wire										w_hcmd_nlb_wr0_en;
wire	[P_SLOT_TAG_WIDTH-1:0]				w_hcmd_nlb_wr0_addr; //slot_modified
wire	[18:0]								w_hcmd_nlb_wr0_data;
wire										w_hcmd_nlb_wr0_rdy_n;

wire										w_hcmd_slot_rdy;
wire	[P_SLOT_TAG_WIDTH-1:0]				w_hcmd_slot_tag; //slot_modified
wire										w_hcmd_slot_alloc_en;

wire										w_hcmd_slot_free_en;
wire	[P_SLOT_TAG_WIDTH-1:0]				w_hcmd_slot_invalid_tag; //slot_modified

wire	[7:0]								w_admin_sq_head_ptr;
wire	[7:0]								w_io_sq1_head_ptr;
wire	[7:0]								w_io_sq2_head_ptr;
wire	[7:0]								w_io_sq3_head_ptr;
wire	[7:0]								w_io_sq4_head_ptr;
wire	[7:0]								w_io_sq5_head_ptr;
wire	[7:0]								w_io_sq6_head_ptr;
wire	[7:0]								w_io_sq7_head_ptr;
wire	[7:0]								w_io_sq8_head_ptr;


pcie_hcmd_table # (
	.P_SLOT_TAG_WIDTH						(P_SLOT_TAG_WIDTH) //slot_modified
)
pcie_hcmd_table_inst0(
	.wr_clk									(pcie_user_clk),

	.wr_en									(w_hcmd_table_wr_en),
	.wr_addr								(w_hcmd_table_wr_addr),
	.wr_data								(w_hcmd_table_wr_data),

	.rd_clk									(cpu_bus_clk),

	.rd_addr								(hcmd_table_rd_addr),
	.rd_data								(hcmd_table_rd_data)
);

pcie_hcmd_table_cid # (
	.P_SLOT_TAG_WIDTH						(P_SLOT_TAG_WIDTH) //slot_modified
)
pcie_hcmd_table_cid_isnt0(
	.clk									(pcie_user_clk),

	.wr_en									(w_hcmd_cid_wr_en),
	.wr_addr								(w_hcmd_cid_wr_addr),
	.wr_data								(w_hcmd_cid_wr_data),

	.rd_addr								(w_hcmd_cid_rd_addr),
	.rd_data								(w_hcmd_cid_rd_data)
);

pcie_hcmd_table_prp # (
	.P_SLOT_TAG_WIDTH						(P_SLOT_TAG_WIDTH) //slot_modified
)
pcie_hcmd_table_prp_isnt0(
	.clk									(pcie_user_clk),

	.wr_en									(w_hcmd_prp_wr_en),
	.wr_addr								(w_hcmd_prp_wr_addr),
	.wr_data								(w_hcmd_prp_wr_data),

	.rd_addr								(hcmd_prp_rd_addr),
	.rd_data								(hcmd_prp_rd_data)
);

pcie_hcmd_nlb # (
	.P_SLOT_TAG_WIDTH						(P_SLOT_TAG_WIDTH) //slot_modified
)
pcie_hcmd_nlb_inst0
(
	.clk									(pcie_user_clk),
	.rst_n									(pcie_user_rst_n),

	.wr0_en									(w_hcmd_nlb_wr0_en),
	.wr0_addr								(w_hcmd_nlb_wr0_addr),
	.wr0_data								(w_hcmd_nlb_wr0_data),
	.wr0_rdy_n								(w_hcmd_nlb_wr0_rdy_n),

	.wr1_en									(hcmd_nlb_wr1_en),
	.wr1_addr								(hcmd_nlb_wr1_addr),
	.wr1_data								(hcmd_nlb_wr1_data),
	.wr1_rdy_n								(hcmd_nlb_wr1_rdy_n),

	.rd_addr								(hcmd_nlb_rd_addr),
	.rd_data								(hcmd_nlb_rd_data)
);

pcie_hcmd_slot_mgt # (
	.P_SLOT_TAG_WIDTH						(P_SLOT_TAG_WIDTH), //slot_modified
	.P_SLOT_WIDTH							(P_SLOT_WIDTH)
)
pcie_hcmd_slot_mgt_inst0
(
	.pcie_user_clk							(pcie_user_clk),
	.pcie_user_rst_n						(pcie_user_rst_n),

	.hcmd_slot_rdy							(w_hcmd_slot_rdy),
	.hcmd_slot_tag							(w_hcmd_slot_tag),
	.hcmd_slot_alloc_en						(w_hcmd_slot_alloc_en),

	.hcmd_slot_free_en						(w_hcmd_slot_free_en),
	.hcmd_slot_invalid_tag					(w_hcmd_slot_invalid_tag)
);

pcie_hcmd_sq # (
	.P_SLOT_TAG_WIDTH						(P_SLOT_TAG_WIDTH), //slot_modified
	.C_PCIE_DATA_WIDTH						(C_PCIE_DATA_WIDTH)
)
pcie_hcmd_sq_inst0(
	.pcie_user_clk							(pcie_user_clk),
	.pcie_user_rst_n						(pcie_user_rst_n),

	.admin_sq_bs_addr						(admin_sq_bs_addr),
	.admin_sq_size							(admin_sq_size),

	.admin_sq_tail_ptr						(admin_sq_tail_ptr),
	.io_sq1_tail_ptr						(io_sq1_tail_ptr),
	.io_sq2_tail_ptr						(io_sq2_tail_ptr),
	.io_sq3_tail_ptr						(io_sq3_tail_ptr),
	.io_sq4_tail_ptr						(io_sq4_tail_ptr),
	.io_sq5_tail_ptr						(io_sq5_tail_ptr),
	.io_sq6_tail_ptr						(io_sq6_tail_ptr),
	.io_sq7_tail_ptr						(io_sq7_tail_ptr),
	.io_sq8_tail_ptr						(io_sq8_tail_ptr),

	.admin_sq_head_ptr						(w_admin_sq_head_ptr),
	.io_sq1_head_ptr						(w_io_sq1_head_ptr),
	.io_sq2_head_ptr						(w_io_sq2_head_ptr),
	.io_sq3_head_ptr						(w_io_sq3_head_ptr),
	.io_sq4_head_ptr						(w_io_sq4_head_ptr),
	.io_sq5_head_ptr						(w_io_sq5_head_ptr),
	.io_sq6_head_ptr						(w_io_sq6_head_ptr),
	.io_sq7_head_ptr						(w_io_sq7_head_ptr),
	.io_sq8_head_ptr						(w_io_sq8_head_ptr),

	.hcmd_slot_rdy							(w_hcmd_slot_rdy),
	.hcmd_slot_tag							(w_hcmd_slot_tag),
	.hcmd_slot_alloc_en						(w_hcmd_slot_alloc_en),

	.cpld_sq_fifo_tag						(cpld_sq_fifo_tag),
	.cpld_sq_fifo_wr_data					(cpld_sq_fifo_wr_data),
	.cpld_sq_fifo_wr_en						(cpld_sq_fifo_wr_en),
	.cpld_sq_fifo_tag_last					(cpld_sq_fifo_tag_last),

	.tx_mrd_req								(tx_mrd_req),
	.tx_mrd_tag								(tx_mrd_tag),
	.tx_mrd_len								(tx_mrd_len),
	.tx_mrd_addr							(tx_mrd_addr),
	.tx_mrd_req_ack							(tx_mrd_req_ack),

	.hcmd_table_wr_en						(w_hcmd_table_wr_en),
	.hcmd_table_wr_addr						(w_hcmd_table_wr_addr),
	.hcmd_table_wr_data						(w_hcmd_table_wr_data),

	.hcmd_cid_wr_en							(w_hcmd_cid_wr_en),
	.hcmd_cid_wr_addr						(w_hcmd_cid_wr_addr),
	.hcmd_cid_wr_data						(w_hcmd_cid_wr_data),

	.hcmd_prp_wr_en							(w_hcmd_prp_wr_en),
	.hcmd_prp_wr_addr						(w_hcmd_prp_wr_addr),
	.hcmd_prp_wr_data						(w_hcmd_prp_wr_data),

	.hcmd_nlb_wr0_en						(w_hcmd_nlb_wr0_en),
	.hcmd_nlb_wr0_addr						(w_hcmd_nlb_wr0_addr),
	.hcmd_nlb_wr0_data						(w_hcmd_nlb_wr0_data),
	.hcmd_nlb_wr0_rdy_n						(w_hcmd_nlb_wr0_rdy_n),

	.cpu_bus_clk							(cpu_bus_clk),
	.cpu_bus_rst_n							(cpu_bus_rst_n),

	.sq_rst_n								(sq_rst_n),
	.sq_valid								(sq_valid),
	.io_sq1_size							(io_sq1_size),
	.io_sq2_size							(io_sq2_size),
	.io_sq3_size							(io_sq3_size),
	.io_sq4_size							(io_sq4_size),
	.io_sq5_size							(io_sq5_size),
	.io_sq6_size							(io_sq6_size),
	.io_sq7_size							(io_sq7_size),
	.io_sq8_size							(io_sq8_size),
	.io_sq1_bs_addr							(io_sq1_bs_addr),
	.io_sq2_bs_addr							(io_sq2_bs_addr),
	.io_sq3_bs_addr							(io_sq3_bs_addr),
	.io_sq4_bs_addr							(io_sq4_bs_addr),
	.io_sq5_bs_addr							(io_sq5_bs_addr),
	.io_sq6_bs_addr							(io_sq6_bs_addr),
	.io_sq7_bs_addr							(io_sq7_bs_addr),
	.io_sq8_bs_addr							(io_sq8_bs_addr),

	.hcmd_sq_rd_en							(hcmd_sq_rd_en),
	.hcmd_sq_rd_data						(hcmd_sq_rd_data),
	.hcmd_sq_empty_n						(hcmd_sq_empty_n)
);

pcie_hcmd_cq # (
	.P_SLOT_TAG_WIDTH						(P_SLOT_TAG_WIDTH), //slot_modified
	.C_PCIE_DATA_WIDTH						(C_PCIE_DATA_WIDTH)
)
pcie_hcmd_cq_inst0(
	.pcie_user_clk							(pcie_user_clk),
	.pcie_user_rst_n						(pcie_user_rst_n),

	.hcmd_cid_rd_addr						(w_hcmd_cid_rd_addr),
	.hcmd_cid_rd_data						(w_hcmd_cid_rd_data),

	.admin_cq_bs_addr						(admin_cq_bs_addr),
	.admin_cq_size							(admin_cq_size),

	.admin_cq_tail_ptr						(admin_cq_tail_ptr),
	.io_cq1_tail_ptr						(io_cq1_tail_ptr),
	.io_cq2_tail_ptr						(io_cq2_tail_ptr),
	.io_cq3_tail_ptr						(io_cq3_tail_ptr),
	.io_cq4_tail_ptr						(io_cq4_tail_ptr),
	.io_cq5_tail_ptr						(io_cq5_tail_ptr),
	.io_cq6_tail_ptr						(io_cq6_tail_ptr),
	.io_cq7_tail_ptr						(io_cq7_tail_ptr),
	.io_cq8_tail_ptr						(io_cq8_tail_ptr),

	.admin_sq_head_ptr						(w_admin_sq_head_ptr),
	.io_sq1_head_ptr						(w_io_sq1_head_ptr),
	.io_sq2_head_ptr						(w_io_sq2_head_ptr),
	.io_sq3_head_ptr						(w_io_sq3_head_ptr),
	.io_sq4_head_ptr						(w_io_sq4_head_ptr),
	.io_sq5_head_ptr						(w_io_sq5_head_ptr),
	.io_sq6_head_ptr						(w_io_sq6_head_ptr),
	.io_sq7_head_ptr						(w_io_sq7_head_ptr),
	.io_sq8_head_ptr						(w_io_sq8_head_ptr),

	.hcmd_slot_free_en						(w_hcmd_slot_free_en),
	.hcmd_slot_invalid_tag					(w_hcmd_slot_invalid_tag),

	.tx_cq_mwr_req							(tx_cq_mwr_req),
	.tx_cq_mwr_tag							(tx_cq_mwr_tag),
	.tx_cq_mwr_len							(tx_cq_mwr_len),
	.tx_cq_mwr_addr							(tx_cq_mwr_addr),
	.tx_cq_mwr_req_ack						(tx_cq_mwr_req_ack),
	.tx_cq_mwr_rd_en						(tx_cq_mwr_rd_en),
	.tx_cq_mwr_rd_data						(tx_cq_mwr_rd_data),
	.tx_cq_mwr_data_last					(tx_cq_mwr_data_last),

	.hcmd_cq_wr0_en							(hcmd_cq_wr0_en),
	.hcmd_cq_wr0_data0						(hcmd_cq_wr0_data0),
	.hcmd_cq_wr0_data1						(hcmd_cq_wr0_data1),
	.hcmd_cq_wr0_rdy_n						(hcmd_cq_wr0_rdy_n),

	.cpu_bus_clk							(cpu_bus_clk),
	.cpu_bus_rst_n							(cpu_bus_rst_n),

	.io_sq1_cq_vec							(io_sq1_cq_vec),
	.io_sq2_cq_vec							(io_sq2_cq_vec),
	.io_sq3_cq_vec							(io_sq3_cq_vec),
	.io_sq4_cq_vec							(io_sq4_cq_vec),
	.io_sq5_cq_vec							(io_sq5_cq_vec),
	.io_sq6_cq_vec							(io_sq6_cq_vec),
	.io_sq7_cq_vec							(io_sq7_cq_vec),
	.io_sq8_cq_vec							(io_sq8_cq_vec),

	.sq_valid								(sq_valid),
	.cq_rst_n								(cq_rst_n),
	.cq_valid								(cq_valid),
	.io_cq1_size							(io_cq1_size),
	.io_cq2_size							(io_cq2_size),
	.io_cq3_size							(io_cq3_size),
	.io_cq4_size							(io_cq4_size),
	.io_cq5_size							(io_cq5_size),
	.io_cq6_size							(io_cq6_size),
	.io_cq7_size							(io_cq7_size),
	.io_cq8_size							(io_cq8_size),
	.io_cq1_bs_addr							(io_cq1_bs_addr),
	.io_cq2_bs_addr							(io_cq2_bs_addr),
	.io_cq3_bs_addr							(io_cq3_bs_addr),
	.io_cq4_bs_addr							(io_cq4_bs_addr),
	.io_cq5_bs_addr							(io_cq5_bs_addr),
	.io_cq6_bs_addr							(io_cq6_bs_addr),
	.io_cq7_bs_addr							(io_cq7_bs_addr),
	.io_cq8_bs_addr							(io_cq8_bs_addr),

	.hcmd_cq_wr1_en							(hcmd_cq_wr1_en),
	.hcmd_cq_wr1_data0						(hcmd_cq_wr1_data0),
	.hcmd_cq_wr1_data1						(hcmd_cq_wr1_data1),
	.hcmd_cq_wr1_rdy_n						(hcmd_cq_wr1_rdy_n)
);

endmodule
