


`timescale 1ns / 1ps

module pcie_hcmd_sq # (
	parameter	C_PCIE_DATA_WIDTH			= 512,
	parameter	C_PCIE_ADDR_WIDTH			= 48, //modified
	parameter 	P_SLOT_TAG_WIDTH			= 10, //slot_modified
	parameter	P_FIFO_DATA_WIDTH			= 128
)
(
	input									pcie_user_clk,
	input									pcie_user_rst_n,
	
	input	[C_PCIE_ADDR_WIDTH-1:2]			admin_sq_bs_addr,
	input	[7:0]							admin_sq_size,

	input	[7:0]							admin_sq_tail_ptr,
	input	[7:0]							io_sq1_tail_ptr,
	input	[7:0]							io_sq2_tail_ptr,
	input	[7:0]							io_sq3_tail_ptr,
	input	[7:0]							io_sq4_tail_ptr,
	input	[7:0]							io_sq5_tail_ptr,
	input	[7:0]							io_sq6_tail_ptr,
	input	[7:0]							io_sq7_tail_ptr,
	input	[7:0]							io_sq8_tail_ptr,

	output	[7:0]							admin_sq_head_ptr,
	output	[7:0]							io_sq1_head_ptr,
	output	[7:0]							io_sq2_head_ptr,
	output	[7:0]							io_sq3_head_ptr,
	output	[7:0]							io_sq4_head_ptr,
	output	[7:0]							io_sq5_head_ptr,
	output	[7:0]							io_sq6_head_ptr,
	output	[7:0]							io_sq7_head_ptr,
	output	[7:0]							io_sq8_head_ptr,

	input									hcmd_slot_rdy,
	input	[P_SLOT_TAG_WIDTH-1:0]			hcmd_slot_tag, //slot_modified
	output									hcmd_slot_alloc_en,

	input	[7:0]							cpld_sq_fifo_tag,
	input	[C_PCIE_DATA_WIDTH-1:0]			cpld_sq_fifo_wr_data,
	input									cpld_sq_fifo_wr_en,
	input									cpld_sq_fifo_tag_last,

	output									tx_mrd_req,
	output	[7:0]							tx_mrd_tag,
	output	[12:2]							tx_mrd_len,
	output	[C_PCIE_ADDR_WIDTH-1:2]			tx_mrd_addr,
	input									tx_mrd_req_ack,

	output									hcmd_table_wr_en,
	output	[(P_SLOT_TAG_WIDTH+2)-1:0]		hcmd_table_wr_addr, //slot_modified
	output	[P_FIFO_DATA_WIDTH-1:0]			hcmd_table_wr_data, 

	output									hcmd_cid_wr_en,
	output	[P_SLOT_TAG_WIDTH-1:0]			hcmd_cid_wr_addr, //slot_modified
	output	[19:0]							hcmd_cid_wr_data,

	output									hcmd_prp_wr_en,
	output	[(P_SLOT_TAG_WIDTH+1)-1:0]		hcmd_prp_wr_addr, //slot_modified
	output	[53:0]							hcmd_prp_wr_data, //modified

	output									hcmd_nlb_wr0_en,
	output	[P_SLOT_TAG_WIDTH-1:0]			hcmd_nlb_wr0_addr, //slot_modified
	output	[18:0]							hcmd_nlb_wr0_data,
	input									hcmd_nlb_wr0_rdy_n,

	input									cpu_bus_clk,
	input									cpu_bus_rst_n,

	input	[8:0]							sq_rst_n,
	input	[8:0]							sq_valid,
	input	[7:0]							io_sq1_size,
	input	[7:0]							io_sq2_size,
	input	[7:0]							io_sq3_size,
	input	[7:0]							io_sq4_size,
	input	[7:0]							io_sq5_size,
	input	[7:0]							io_sq6_size,
	input	[7:0]							io_sq7_size,
	input	[7:0]							io_sq8_size,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq1_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq2_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq3_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq4_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq5_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq6_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq7_bs_addr,
	input	[C_PCIE_ADDR_WIDTH-1:2]			io_sq8_bs_addr,

	input									hcmd_sq_rd_en,
	output	[(P_SLOT_TAG_WIDTH+12)-1:0]		hcmd_sq_rd_data, //slot_modified
	output									hcmd_sq_empty_n
);

wire										w_arb_sq_rdy;
wire	[3:0]								w_sq_qid;
wire	[C_PCIE_ADDR_WIDTH-1:2]				w_hcmd_pcie_addr;
wire										w_sq_hcmd_ack;

wire										w_hcmd_sq_wr_en;
wire	[(P_SLOT_TAG_WIDTH+12)-1:0]			w_hcmd_sq_wr_data; //slot_modified
wire										w_hcmd_sq_full_n;

wire										w_pcie_sq_cmd_fifo_wr_en;
wire	[(P_SLOT_TAG_WIDTH+4)-1:0]			w_pcie_sq_cmd_fifo_wr_data; //slot_modified
wire										w_pcie_sq_cmd_fifo_full_n;

wire										w_pcie_sq_cmd_fifo_rd_en;
wire	[(P_SLOT_TAG_WIDTH+4)-1:0]			w_pcie_sq_cmd_fifo_rd_data; //slot_modified
wire										w_pcie_sq_cmd_fifo_empty_n;

wire										w_pcie_sq_rx_tag_alloc;
wire	[7:0]								w_pcie_sq_rx_alloc_tag;
wire									w_pcie_sq_rx_tag_alloc_len;
wire										w_pcie_sq_rx_tag_full_n;

wire										w_pcie_sq_rx_fifo_wr_en;
wire	[3:0]								w_pcie_sq_rx_fifo_wr_addr;
wire	[C_PCIE_DATA_WIDTH-1:0]				w_pcie_sq_rx_fifo_wr_data;
wire	[4:0]								w_pcie_sq_rx_fifo_rear_full_addr;
wire	[4:0]								w_pcie_sq_rx_fifo_rear_addr;
wire										w_pcie_sq_rx_fifo_full_n;

wire										w_pcie_sq_rx_fifo_rd_en;
wire	[C_PCIE_DATA_WIDTH-1:0]				w_pcie_sq_rx_fifo_rd_data;
wire										w_pcie_sq_rx_fifo_free_en;
wire									w_pcie_sq_rx_fifo_free_len;
wire										w_pcie_sq_rx_fifo_empty_n;


pcie_hcmd_sq_fifo # (
	.P_SLOT_TAG_WIDTH						(P_SLOT_TAG_WIDTH) //slot_modified
)
pcie_hcmd_sq_fifo_inst0(
	.wr_clk									(pcie_user_clk),
	.wr_rst_n								(pcie_user_rst_n),

	.wr_en									(w_hcmd_sq_wr_en),
	.wr_data								(w_hcmd_sq_wr_data),
	.full_n									(w_hcmd_sq_full_n),

	.rd_clk									(cpu_bus_clk),
	.rd_rst_n								(pcie_user_rst_n),

	.rd_en									(hcmd_sq_rd_en),
	.rd_data								(hcmd_sq_rd_data),
	.empty_n								(hcmd_sq_empty_n)
);

pcie_sq_cmd_fifo # (
	.P_SLOT_TAG_WIDTH						(P_SLOT_TAG_WIDTH) //slot_modified
)
pcie_sq_cmd_fifo_inst0
(
	.clk									(pcie_user_clk),
	.rst_n									(pcie_user_rst_n),

	.wr_en									(w_pcie_sq_cmd_fifo_wr_en),
	.wr_data								(w_pcie_sq_cmd_fifo_wr_data),
	.full_n									(w_pcie_sq_cmd_fifo_full_n),

	.rd_en									(w_pcie_sq_cmd_fifo_rd_en),
	.rd_data								(w_pcie_sq_cmd_fifo_rd_data),
	.empty_n								(w_pcie_sq_cmd_fifo_empty_n)
);

pcie_sq_rx_fifo
pcie_sq_rx_fifo_inst0
(
	.clk									(pcie_user_clk),
	.rst_n									(pcie_user_rst_n),

	.wr_en									(w_pcie_sq_rx_fifo_wr_en),
	.wr_addr								(w_pcie_sq_rx_fifo_wr_addr),
	.wr_data								(w_pcie_sq_rx_fifo_wr_data),
	.rear_full_addr							(w_pcie_sq_rx_fifo_rear_full_addr),
	.rear_addr								(w_pcie_sq_rx_fifo_rear_addr),
	.alloc_len								(w_pcie_sq_rx_tag_alloc_len),
	.full_n									(w_pcie_sq_rx_fifo_full_n),

	.rd_en									(w_pcie_sq_rx_fifo_rd_en),
	.rd_data								(w_pcie_sq_rx_fifo_rd_data),
	.free_en								(w_pcie_sq_rx_fifo_free_en),
	.free_len								(w_pcie_sq_rx_fifo_free_len),
	.empty_n								(w_pcie_sq_rx_fifo_empty_n)
);

pcie_sq_rx_tag
pcie_sq_rx_tag_inst0
(
	.pcie_user_clk							(pcie_user_clk),
	.pcie_user_rst_n						(pcie_user_rst_n),

	.pcie_tag_alloc							(w_pcie_sq_rx_tag_alloc),
	.pcie_alloc_tag							(w_pcie_sq_rx_alloc_tag),
	.pcie_tag_alloc_len						(w_pcie_sq_rx_tag_alloc_len),
	.pcie_tag_full_n						(w_pcie_sq_rx_tag_full_n),

	.cpld_fifo_tag							(cpld_sq_fifo_tag),
	.cpld_fifo_wr_data						(cpld_sq_fifo_wr_data),
	.cpld_fifo_wr_en						(cpld_sq_fifo_wr_en),
	.cpld_fifo_tag_last						(cpld_sq_fifo_tag_last),

	.fifo_wr_en								(w_pcie_sq_rx_fifo_wr_en),
	.fifo_wr_addr							(w_pcie_sq_rx_fifo_wr_addr),
	.fifo_wr_data							(w_pcie_sq_rx_fifo_wr_data),
	.rear_full_addr							(w_pcie_sq_rx_fifo_rear_full_addr),
	.rear_addr								(w_pcie_sq_rx_fifo_rear_addr)
);

pcie_hcmd_sq_arb
pcie_hcmd_sq_arb_inst0
(
	.pcie_user_clk							(pcie_user_clk),
	.pcie_user_rst_n						(pcie_user_rst_n),

	.sq_rst_n								(sq_rst_n),
	.sq_valid								(sq_valid),
	.admin_sq_size							(admin_sq_size),
	.io_sq1_size							(io_sq1_size),
	.io_sq2_size							(io_sq2_size),
	.io_sq3_size							(io_sq3_size),
	.io_sq4_size							(io_sq4_size),
	.io_sq5_size							(io_sq5_size),
	.io_sq6_size							(io_sq6_size),
	.io_sq7_size							(io_sq7_size),
	.io_sq8_size							(io_sq8_size),
	.admin_sq_bs_addr						(admin_sq_bs_addr),
	.io_sq1_bs_addr							(io_sq1_bs_addr),
	.io_sq2_bs_addr							(io_sq2_bs_addr),
	.io_sq3_bs_addr							(io_sq3_bs_addr),
	.io_sq4_bs_addr							(io_sq4_bs_addr),
	.io_sq5_bs_addr							(io_sq5_bs_addr),
	.io_sq6_bs_addr							(io_sq6_bs_addr),
	.io_sq7_bs_addr							(io_sq7_bs_addr),
	.io_sq8_bs_addr							(io_sq8_bs_addr),

	.admin_sq_tail_ptr						(admin_sq_tail_ptr),
	.io_sq1_tail_ptr						(io_sq1_tail_ptr),
	.io_sq2_tail_ptr						(io_sq2_tail_ptr),
	.io_sq3_tail_ptr						(io_sq3_tail_ptr),
	.io_sq4_tail_ptr						(io_sq4_tail_ptr),
	.io_sq5_tail_ptr						(io_sq5_tail_ptr),
	.io_sq6_tail_ptr						(io_sq6_tail_ptr),
	.io_sq7_tail_ptr						(io_sq7_tail_ptr),
	.io_sq8_tail_ptr						(io_sq8_tail_ptr),

	.arb_sq_rdy								(w_arb_sq_rdy),
	.sq_qid									(w_sq_qid),
	.hcmd_pcie_addr							(w_hcmd_pcie_addr),
	.sq_hcmd_ack							(w_sq_hcmd_ack)
);

pcie_hcmd_sq_req # (
	.P_SLOT_TAG_WIDTH						(P_SLOT_TAG_WIDTH), //slot_modified
	.C_PCIE_DATA_WIDTH						(C_PCIE_DATA_WIDTH)
)
pcie_hcmd_sq_req_inst0(
	.pcie_user_clk							(pcie_user_clk),
	.pcie_user_rst_n						(pcie_user_rst_n),

	.arb_sq_rdy								(w_arb_sq_rdy),
	.sq_qid									(w_sq_qid),
	.hcmd_pcie_addr							(w_hcmd_pcie_addr),
	.sq_hcmd_ack							(w_sq_hcmd_ack),

	.hcmd_slot_rdy							(hcmd_slot_rdy),
	.hcmd_slot_tag							(hcmd_slot_tag),
	.hcmd_slot_alloc_en						(hcmd_slot_alloc_en),

	.pcie_sq_cmd_fifo_wr_en					(w_pcie_sq_cmd_fifo_wr_en),
	.pcie_sq_cmd_fifo_wr_data				(w_pcie_sq_cmd_fifo_wr_data),
	.pcie_sq_cmd_fifo_full_n				(w_pcie_sq_cmd_fifo_full_n),

	.pcie_sq_rx_tag_alloc					(w_pcie_sq_rx_tag_alloc),
	.pcie_sq_rx_alloc_tag					(w_pcie_sq_rx_alloc_tag),
	.pcie_sq_rx_tag_alloc_len				(w_pcie_sq_rx_tag_alloc_len),
	.pcie_sq_rx_tag_full_n					(w_pcie_sq_rx_tag_full_n),
	.pcie_sq_rx_fifo_full_n					(w_pcie_sq_rx_fifo_full_n),

	.tx_mrd_req								(tx_mrd_req),
	.tx_mrd_tag								(tx_mrd_tag),
	.tx_mrd_len								(tx_mrd_len),
	.tx_mrd_addr							(tx_mrd_addr),
	.tx_mrd_req_ack							(tx_mrd_req_ack)
);


pcie_hcmd_sq_recv # (
	.P_SLOT_TAG_WIDTH						(P_SLOT_TAG_WIDTH) //slot_modified
)
pcie_hcmd_sq_recv_inst0
(
	.pcie_user_clk							(pcie_user_clk),
	.pcie_user_rst_n						(pcie_user_rst_n),
	
	.pcie_sq_cmd_fifo_rd_en					(w_pcie_sq_cmd_fifo_rd_en),
	.pcie_sq_cmd_fifo_rd_data				(w_pcie_sq_cmd_fifo_rd_data),
	.pcie_sq_cmd_fifo_empty_n				(w_pcie_sq_cmd_fifo_empty_n),

	.pcie_sq_rx_fifo_rd_en					(w_pcie_sq_rx_fifo_rd_en),
	.pcie_sq_rx_fifo_rd_data				(w_pcie_sq_rx_fifo_rd_data),
	.pcie_sq_rx_fifo_free_en				(w_pcie_sq_rx_fifo_free_en),
	.pcie_sq_rx_fifo_free_len				(w_pcie_sq_rx_fifo_free_len),
	.pcie_sq_rx_fifo_empty_n				(w_pcie_sq_rx_fifo_empty_n),

	.hcmd_table_wr_en						(hcmd_table_wr_en),
	.hcmd_table_wr_addr						(hcmd_table_wr_addr),
	.hcmd_table_wr_data						(hcmd_table_wr_data),

	.hcmd_cid_wr_en							(hcmd_cid_wr_en),
	.hcmd_cid_wr_addr						(hcmd_cid_wr_addr),
	.hcmd_cid_wr_data						(hcmd_cid_wr_data),

	.hcmd_prp_wr_en							(hcmd_prp_wr_en),
	.hcmd_prp_wr_addr						(hcmd_prp_wr_addr),
	.hcmd_prp_wr_data						(hcmd_prp_wr_data),

	.hcmd_nlb_wr0_en						(hcmd_nlb_wr0_en),
	.hcmd_nlb_wr0_addr						(hcmd_nlb_wr0_addr),
	.hcmd_nlb_wr0_data						(hcmd_nlb_wr0_data),
	.hcmd_nlb_wr0_rdy_n						(hcmd_nlb_wr0_rdy_n),

	.hcmd_sq_wr_en							(w_hcmd_sq_wr_en),
	.hcmd_sq_wr_data						(w_hcmd_sq_wr_data),
	.hcmd_sq_full_n							(w_hcmd_sq_full_n),

	.sq_rst_n								(sq_rst_n),
	.admin_sq_size							(admin_sq_size),
	.io_sq1_size							(io_sq1_size),
	.io_sq2_size							(io_sq2_size),
	.io_sq3_size							(io_sq3_size),
	.io_sq4_size							(io_sq4_size),
	.io_sq5_size							(io_sq5_size),
	.io_sq6_size							(io_sq6_size),
	.io_sq7_size							(io_sq7_size),
	.io_sq8_size							(io_sq8_size),

	.admin_sq_head_ptr						(admin_sq_head_ptr),
	.io_sq1_head_ptr						(io_sq1_head_ptr),
	.io_sq2_head_ptr						(io_sq2_head_ptr),
	.io_sq3_head_ptr						(io_sq3_head_ptr),
	.io_sq4_head_ptr						(io_sq4_head_ptr),
	.io_sq5_head_ptr						(io_sq5_head_ptr),
	.io_sq6_head_ptr						(io_sq6_head_ptr),
	.io_sq7_head_ptr						(io_sq7_head_ptr),
	.io_sq8_head_ptr						(io_sq8_head_ptr)
);

endmodule
