


`timescale 1ns / 1ps

`include	"def_axi.vh"

 module m_axi_write # (
	parameter 	P_SLOT_TAG_WIDTH			=  10, //slot_modified
	parameter	C_M_AXI_ADDR_WIDTH			= 32,
	parameter	C_M_AXI_DATA_WIDTH			= 64,
	parameter	C_M_AXI_ID_WIDTH			= 1,
	parameter	C_M_AXI_AWUSER_WIDTH		= 1,
	parameter	C_M_AXI_WUSER_WIDTH			= 1,
	parameter	C_M_AXI_BUSER_WIDTH			= 1
)
(

////////////////////////////////////////////////////////////////
//AXI4 master write channel signal
 	input									m_axi_aclk,
 	input									m_axi_aresetn,

	// Write address channel
 	output	[C_M_AXI_ID_WIDTH-1:0]			m_axi_awid,
 	output	[C_M_AXI_ADDR_WIDTH-1:0]		m_axi_awaddr,
 	output	[7:0]							m_axi_awlen,
 	output	[2:0]							m_axi_awsize,
 	output	[1:0]							m_axi_awburst,
 	output	[1:0]							m_axi_awlock,
	 output	[3:0]							m_axi_awcache,
	 output	[2:0]							m_axi_awprot,
	 output	[3:0]							m_axi_awregion,
	 output	[3:0]							m_axi_awqos,
	 output	[C_M_AXI_AWUSER_WIDTH-1:0]		m_axi_awuser,
	 output									m_axi_awvalid,
	 input									m_axi_awready,

// Write data channel
 	output	[C_M_AXI_ID_WIDTH-1:0]			m_axi_wid,
 	output	[C_M_AXI_DATA_WIDTH-1:0]		m_axi_wdata,
	 output	[(C_M_AXI_DATA_WIDTH/8)-1:0]	m_axi_wstrb,
	 output									m_axi_wlast,
 	output	[C_M_AXI_WUSER_WIDTH-1:0]		m_axi_wuser,
 	output									m_axi_wvalid,
 	input									m_axi_wready,

// Write response channel
 	input	[C_M_AXI_ID_WIDTH-1:0]			m_axi_bid,
 	input	[1:0]							m_axi_bresp,
 	input									m_axi_bvalid,
 	input	[C_M_AXI_BUSER_WIDTH-1:0]		m_axi_buser,
	 output									m_axi_bready,

 	output									m_axi_bresp_err,

 	output									dev_rx_cmd_rd_en,
 	input	[29:0]							dev_rx_cmd_rd_data,
 	input									dev_rx_cmd_empty_n,

 	output									pcie_rx_fifo_rd_en,
 	input	[C_M_AXI_DATA_WIDTH-1:0]		pcie_rx_fifo_rd_data,
 	output									pcie_rx_fifo_free_en,
 	output	[10:6]							pcie_rx_fifo_free_len,
 	input									pcie_rx_fifo_empty_n,

 	output									dma_rx_done_wr_en,
	 output	[(P_SLOT_TAG_WIDTH+15)-1:0]		dma_rx_done_wr_data,
	 input									dma_rx_done_wr_rdy_n
);

localparam	LP_AW_DELAY						= 7;

localparam	S_AW_IDLE						= 11'b00000000001;
localparam	S_AW_CMD_0						= 11'b00000000010;
localparam	S_AW_CMD_1						= 11'b00000000100;
localparam	S_AW_WAIT_EMPTY_N				= 11'b00000001000;
localparam	S_AW_REQ						= 11'b00000010000;
localparam	S_AW_WAIT						= 11'b00000100000;
localparam	S_AW_W_REQ						= 11'b00001000000;
localparam	S_AW_DONE						= 11'b00010000000;
localparam	S_AW_DELAY						= 11'b00100000000;
localparam	S_AW_DMA_DONE_WR_WAIT			= 11'b01000000000;
localparam	S_AW_DMA_DONE_WR				= 11'b10000000000;

     reg		[10:0]								cur_aw_state;
     reg		[10:0]								next_aw_state;
    
    localparam	S_W_IDLE						= 4'b0001;
    localparam	S_W_DATA						= 4'b0010;
    localparam	S_W_READY_WAIT					= 4'b0100;
    localparam	S_W_DATA_LAST					= 4'b1000;
    
    reg		[4:0]								cur_w_state;
     reg		[4:0]								next_w_state;
    
     reg											r_dma_cmd_type;
     reg											r_dma_cmd_auto_cpl;
     reg											r_dma_done_check;
     reg		[P_SLOT_TAG_WIDTH-1:0]				r_hcmd_slot_tag; //slot_modified
     reg		[31:2]								r_dev_addr;
     reg		[31:2]								r_dev_addr_backup;     
     reg		[12:2]								r_dev_dma_len;
     reg		[12:2]								r_dev_dma_orig_len;
     reg		[10:2]								r_dev_cur_len;
     reg		[10:2]								r_wr_data_cnt;
     reg		[4:0]								r_aw_delay;
       
     reg		[10:2]								r_m_axi_awlen;
     reg											r_m_axi_awvalid;
     reg		[C_M_AXI_DATA_WIDTH-1:0]			r_m_axi_wdata;
     reg											r_m_axi_wlast;
     reg											r_m_axi_wvalid;
     reg											r_m_axi_wdata_sel;
    
     reg											r_m_axi_bvalid;
    //reg											r_m_axi_bvalid_d1;
    //wire										w_m_axi_bvalid;
     reg		[C_M_AXI_ID_WIDTH-1:0]				r_m_axi_bid;
    reg		[1:0]								r_m_axi_bresp;
     reg											r_m_axi_bresp_err;
     reg											r_m_axi_bresp_err_d1;
     reg											r_m_axi_bresp_err_d2;
    
     reg		[2:0]								r_axi_aw_req_gnt;
     reg											r_axi_aw_req;
     wire										w_axi_aw_req_gnt;
     reg											r_axi_wr_req;
     reg											r_axi_wr_rdy;
    
     reg											r_dev_rx_cmd_rd_en;
     reg											r_pcie_rx_fifo_rd_en;
     reg		[C_M_AXI_DATA_WIDTH-1:0]			r_pcie_rx_fifo_rd_data;
     reg		[C_M_AXI_DATA_WIDTH-1:0]			r_pcie_rx_fifo_rd_data_d1;
     reg											r_pcie_rx_fifo_free_en;
    
     reg											r_dma_rx_done_wr_en;

 	reg			[2:0]                               r_wr_count;
	reg                                             r_dummy_write;
	reg			[10:6]								r_pcie_rx_fifo_free_len;
	 reg											r_2nd_dma;
     wire	[63:0]								w_one_padding;

assign w_one_padding = 64'hFFFF_FFFF_FFFF_FFFF;

assign m_axi_awid = 0;
assign m_axi_awaddr = {r_dev_addr, 2'b0};
assign m_axi_awlen = r_m_axi_awlen[10:3];
assign m_axi_awsize = `D_AXSIZE_008_BYTES;
assign m_axi_awburst = `D_AXBURST_INCR;
assign m_axi_awlock = `D_AXLOCK_NORMAL;
assign m_axi_awcache = `D_AXCACHE_NON_CACHE;
assign m_axi_awprot = `D_AXPROT_SECURE;
assign m_axi_awregion = 0;
assign m_axi_awqos = 0;
assign m_axi_awuser = 0;
assign m_axi_awvalid = r_m_axi_awvalid;

assign m_axi_wid = 0;
assign m_axi_wdata = r_m_axi_wdata;
assign m_axi_wstrb = w_one_padding[(C_M_AXI_DATA_WIDTH/8)-1:0];
assign m_axi_wlast = r_m_axi_wlast;
assign m_axi_wuser = 0;
assign m_axi_wvalid = r_m_axi_wvalid;

assign m_axi_bready = 1;
assign m_axi_bresp_err = r_m_axi_bresp_err_d2;

assign dev_rx_cmd_rd_en = r_dev_rx_cmd_rd_en;
assign pcie_rx_fifo_rd_en = r_pcie_rx_fifo_rd_en;
assign pcie_rx_fifo_free_en = r_pcie_rx_fifo_free_en;
assign pcie_rx_fifo_free_len = r_pcie_rx_fifo_free_len;

assign dma_rx_done_wr_en = r_dma_rx_done_wr_en;
assign dma_rx_done_wr_data = {r_dma_cmd_auto_cpl, r_dma_cmd_type, r_dma_done_check, 1'b0, r_hcmd_slot_tag, r_dev_dma_orig_len};


always @ (posedge m_axi_aclk or negedge m_axi_aresetn)
begin
	if(m_axi_aresetn == 0)
		cur_aw_state <= S_AW_IDLE;
	else
		cur_aw_state <= next_aw_state;
end

always @ (*)
begin
	case(cur_aw_state)
		S_AW_IDLE: begin
			if(dev_rx_cmd_empty_n == 1)
				next_aw_state <= S_AW_CMD_0;
			else
				next_aw_state <= S_AW_IDLE;
		end
		S_AW_CMD_0: begin
			next_aw_state <= S_AW_CMD_1;
		end
		S_AW_CMD_1: begin
			next_aw_state <= S_AW_WAIT_EMPTY_N;
		end
		S_AW_WAIT_EMPTY_N: begin
			if(pcie_rx_fifo_empty_n == 1 && w_axi_aw_req_gnt == 1)
				next_aw_state <= S_AW_REQ;
			else
				next_aw_state <= S_AW_WAIT_EMPTY_N;
		end
		S_AW_REQ: begin
			if(m_axi_awready == 1)
				next_aw_state <= S_AW_W_REQ;
			else
				next_aw_state <= S_AW_WAIT;
		end
		S_AW_WAIT: begin
			if(m_axi_awready == 1)
				next_aw_state <= S_AW_W_REQ;
			else
				next_aw_state <= S_AW_WAIT;
		end
		S_AW_W_REQ: begin
			if(r_axi_wr_rdy == 1)
				next_aw_state <= S_AW_DONE;
			else
				next_aw_state <= S_AW_W_REQ;
		end
		S_AW_DONE: begin
			if(r_dummy_write != 1 && r_dev_dma_len == 0)
				next_aw_state <= S_AW_DMA_DONE_WR_WAIT;
			else
				next_aw_state <= S_AW_DELAY;
		end
		S_AW_DELAY: begin
			if(r_aw_delay == 0)
				next_aw_state <= S_AW_WAIT_EMPTY_N;
			else
				next_aw_state <= S_AW_DELAY;
		end
		S_AW_DMA_DONE_WR_WAIT: begin
			if(dma_rx_done_wr_rdy_n == 1)
				next_aw_state <= S_AW_DMA_DONE_WR_WAIT;
			else
				next_aw_state <= S_AW_DMA_DONE_WR;
		end
		S_AW_DMA_DONE_WR: begin
			next_aw_state <= S_AW_IDLE;
		end
		default: begin
			next_aw_state <= S_AW_IDLE;
		end
	endcase
end

always @ (posedge m_axi_aclk)
begin
	case(cur_aw_state)
		S_AW_IDLE: begin

		end
		S_AW_CMD_0: begin
		    r_dma_cmd_auto_cpl <= dev_rx_cmd_rd_data[P_SLOT_TAG_WIDTH+13]; //slot_modified
			r_dma_cmd_type     <= dev_rx_cmd_rd_data[P_SLOT_TAG_WIDTH+12]; //slot_modified
			r_dma_done_check   <= dev_rx_cmd_rd_data[P_SLOT_TAG_WIDTH+11];
			r_hcmd_slot_tag    <= dev_rx_cmd_rd_data[(P_SLOT_TAG_WIDTH+11)-1:11]; //slot_modified
			r_dev_dma_len      <= {dev_rx_cmd_rd_data[10:2], 2'b0};
			if(dev_rx_cmd_rd_data[9:2] != 0) begin
				if(r_2nd_dma == 0)
					r_2nd_dma <= 1;
				else
					r_2nd_dma <= 0;
			end
			else
				r_2nd_dma <= 0;
		end
		S_AW_CMD_1: begin
			r_dev_dma_orig_len <= r_dev_dma_len;
			if(r_2nd_dma == 1) begin
				if(r_dev_dma_len[5:2] != 0) begin
					r_dev_cur_len[10:2]           <= {5'b0, r_dev_dma_len[5:2]};
					r_pcie_rx_fifo_free_len[10:6] <= 5'b1;
				end
				else if(r_dev_dma_len[12:2] >= 9'h100) begin
					r_dev_cur_len[10:2]           <= 9'h100;
					r_pcie_rx_fifo_free_len[10:6] <= 5'h10;
				end
				else begin
					r_dev_cur_len[10:2]           <= {1'b0, r_dev_dma_len[9:6], 4'b0};
					r_pcie_rx_fifo_free_len[10:6] <= {1'b0, r_dev_dma_len[9:6]};
				end
			end
			else begin
				if(r_dev_dma_len[12:2] >= 9'h100) begin
					r_dev_cur_len[10:2]           <= 9'h100;
					r_pcie_rx_fifo_free_len[10:6] <= 5'h10;
				end
				else if(r_dev_dma_len[9:6] != 0) begin
					r_dev_cur_len[10:2]           <= {1'b0, r_dev_dma_len[9:6], 4'b0};
					r_pcie_rx_fifo_free_len[10:6] <= {1'b0, r_dev_dma_len[9:6]};
				end
				else begin
					r_dev_cur_len[10:2]           <= {5'b0, r_dev_dma_len[5:2]};
					r_pcie_rx_fifo_free_len[10:6] <= 5'b1;
				end
			end

			r_dev_addr        <= {dev_rx_cmd_rd_data[29:2], 2'b0};
			r_dev_addr_backup <= {dev_rx_cmd_rd_data[29:2], 2'b0};

			if(r_dev_dma_len[5:2] != 0)
				r_wr_count   <= 4'h8 - r_dev_dma_len[5:3] - r_dev_dma_len[2];
			else
				r_wr_count   <= 0;			
			r_dummy_write <= 0;
		end
		S_AW_WAIT_EMPTY_N: begin
			if(r_dummy_write == 1)
				r_m_axi_awlen           <= r_wr_count * 2'b10 - 2;
			else
				r_m_axi_awlen <= r_dev_cur_len - 2;
		end
		S_AW_REQ: begin
			if(r_dummy_write == 1)
				r_wr_count    <= 0;
			else
				r_dev_dma_len <= r_dev_dma_len - r_dev_cur_len;
		end
		S_AW_WAIT: begin
 
		end
		S_AW_W_REQ: begin
			if(r_2nd_dma == 1 && r_wr_count != 0)
				r_dummy_write <= 1;
			else if(r_2nd_dma == 0 && r_dev_dma_len == 0 && r_wr_count != 0)
				r_dummy_write <= 1;
			else
				r_dummy_write <= 0;
		    r_dev_addr        <= r_dev_addr_backup;
		end
		S_AW_DONE: begin
			if(r_dummy_write == 1) begin
			    r_dev_addr                    <= 30'h1FFFF000;
				r_pcie_rx_fifo_free_len[10:6] <= 5'b0;
			end
			else begin
				if(r_2nd_dma == 1) begin
					if(r_dev_dma_len[12:2] >= 9'h100) begin
						r_dev_cur_len[10:2]           <= 9'h100;
						r_pcie_rx_fifo_free_len[10:6] <= 5'h10;
					end
					else begin
						r_dev_cur_len[10:2]           <= {1'b0, r_dev_dma_len[9:6], 4'b0};
						r_pcie_rx_fifo_free_len[10:6] <= {1'b0, r_dev_dma_len[9:6]};
					end
				end
				else begin
					if(r_dev_dma_len[12:2] >= 9'h100) begin
						r_dev_cur_len[10:2]           <= 9'h100;
						r_pcie_rx_fifo_free_len[10:6] <= 5'h10;
					end
					else if(r_dev_dma_len[9:6] != 0) begin
						r_dev_cur_len[10:2]           <= {1'b0, r_dev_dma_len[9:6], 4'b0};
						r_pcie_rx_fifo_free_len[10:6] <= {1'b0, r_dev_dma_len[9:6]};
					end
					else begin
						r_dev_cur_len[10:2]           <= {5'b0, r_dev_dma_len[5:2]};
						r_pcie_rx_fifo_free_len[10:6] <= 5'b1;
					end
				end
				r_dev_addr <= r_dev_addr + r_dev_cur_len;
			end
			r_aw_delay <= LP_AW_DELAY;
		end
		S_AW_DELAY: begin
			r_aw_delay <= r_aw_delay - 1;
			if(r_dummy_write != 1)
			    r_dev_addr_backup   <= r_dev_addr;
		end
		S_AW_DMA_DONE_WR_WAIT: begin

		end
		S_AW_DMA_DONE_WR: begin

		end
		default: begin

		end
	endcase
end


always @ (*)
begin
	case(cur_aw_state)
		S_AW_IDLE: begin
			r_dev_rx_cmd_rd_en <= 0;
			r_m_axi_awvalid <= 0;
			r_axi_aw_req <= 0;
			r_axi_wr_req <= 0;
			r_pcie_rx_fifo_free_en <= 0;
			r_dma_rx_done_wr_en <= 0;
		end
		S_AW_CMD_0: begin
			r_dev_rx_cmd_rd_en <= 1;
			r_m_axi_awvalid <= 0;
			r_axi_aw_req <= 0;
			r_axi_wr_req <= 0;
			r_pcie_rx_fifo_free_en <= 0;
			r_dma_rx_done_wr_en <= 0;
		end
		S_AW_CMD_1: begin
			r_dev_rx_cmd_rd_en <= 1;
			r_m_axi_awvalid <= 0;
			r_axi_aw_req <= 0;
			r_axi_wr_req <= 0;
			r_pcie_rx_fifo_free_en <= 0;
			r_dma_rx_done_wr_en <= 0;
		end
		S_AW_WAIT_EMPTY_N: begin
			r_dev_rx_cmd_rd_en <= 0;
			r_m_axi_awvalid <= 0;
			r_axi_aw_req <= 0;
			r_axi_wr_req <= 0;
			r_pcie_rx_fifo_free_en <= 0;
			r_dma_rx_done_wr_en <= 0;
		end
		S_AW_REQ: begin
			r_dev_rx_cmd_rd_en <= 0;
			r_m_axi_awvalid <= 1;
			r_axi_aw_req <= 1;
			r_axi_wr_req <= 0;
			r_pcie_rx_fifo_free_en <= 1;
			r_dma_rx_done_wr_en <= 0;
		end
		S_AW_WAIT: begin
			r_dev_rx_cmd_rd_en <= 0;
			r_m_axi_awvalid <= 1;
			r_axi_aw_req <= 0;
			r_axi_wr_req <= 0;
			r_pcie_rx_fifo_free_en <= 0;
			r_dma_rx_done_wr_en <= 0;
		end
		S_AW_W_REQ: begin
			r_dev_rx_cmd_rd_en <= 0;
			r_m_axi_awvalid <= 0;
			r_axi_aw_req <= 0;
			r_axi_wr_req <= 1;
			r_pcie_rx_fifo_free_en <= 0;
			r_dma_rx_done_wr_en <= 0;
		end
		S_AW_DONE: begin
			r_dev_rx_cmd_rd_en <= 0;
			r_m_axi_awvalid <= 0;
			r_axi_aw_req <= 0;
			r_axi_wr_req <= 0;
			r_pcie_rx_fifo_free_en <= 0;
			r_dma_rx_done_wr_en <= 0;
		end
		S_AW_DELAY: begin
			r_dev_rx_cmd_rd_en <= 0;
			r_m_axi_awvalid <= 0;
			r_axi_aw_req <= 0;
			r_axi_wr_req <= 0;
			r_pcie_rx_fifo_free_en <= 0;
			r_dma_rx_done_wr_en <= 0;
		end
		S_AW_DMA_DONE_WR_WAIT: begin
			r_dev_rx_cmd_rd_en <= 0;
			r_m_axi_awvalid <= 0;
			r_axi_aw_req <= 0;
			r_axi_wr_req <= 0;
			r_pcie_rx_fifo_free_en <= 0;
			r_dma_rx_done_wr_en <= 0;
		end
		S_AW_DMA_DONE_WR: begin
			r_dev_rx_cmd_rd_en <= 0;
			r_m_axi_awvalid <= 0;
			r_axi_aw_req <= 0;
			r_axi_wr_req <= 0;
			r_pcie_rx_fifo_free_en <= 0;
			r_dma_rx_done_wr_en <= 1;
		end
		default: begin
			r_dev_rx_cmd_rd_en <= 0;
			r_m_axi_awvalid <= 0;
			r_axi_aw_req <= 0;
			r_axi_wr_req <= 0;
			r_pcie_rx_fifo_free_en <= 0;
			r_dma_rx_done_wr_en <= 0;
		end
	endcase
end

assign w_axi_aw_req_gnt = r_axi_aw_req_gnt[2];

//assign w_m_axi_bvalid = r_m_axi_bvalid & ~r_m_axi_bvalid_d1;

always @ (posedge m_axi_aclk)
begin
	r_m_axi_bvalid <= m_axi_bvalid;
//	r_m_axi_bvalid_d1 <= r_m_axi_bvalid;
	r_m_axi_bid <= m_axi_bid;
	r_m_axi_bresp <= m_axi_bresp;

	r_m_axi_bresp_err_d1 <= r_m_axi_bresp_err;
	r_m_axi_bresp_err_d2 <= r_m_axi_bresp_err | r_m_axi_bresp_err_d1;
end

always @ (*)
begin
	if(r_m_axi_bvalid == 1 && (r_m_axi_bresp != `D_AXI_RESP_OKAY || r_m_axi_bid != 0))
		r_m_axi_bresp_err <= 1;
	else
		r_m_axi_bresp_err <= 0;
end

always @ (posedge m_axi_aclk or negedge m_axi_aresetn)
begin
	if(m_axi_aresetn == 0) begin
		r_axi_aw_req_gnt <= 3'b110;
	end
	else begin
		case({r_m_axi_bvalid, r_axi_aw_req})
			2'b01: begin
				r_axi_aw_req_gnt <= {r_axi_aw_req_gnt[1:0], r_axi_aw_req_gnt[2]};
			end
			2'b10: begin
				r_axi_aw_req_gnt <= {r_axi_aw_req_gnt[0], r_axi_aw_req_gnt[2:1]};
			end
			default: begin

			end
		endcase
	end
end

always @ (posedge m_axi_aclk or negedge m_axi_aresetn)
begin
	if(m_axi_aresetn == 0)
		cur_w_state <= S_W_IDLE;
	else
		cur_w_state <= next_w_state;
end

always @ (*)
begin
	case(cur_w_state)
		S_W_IDLE: begin
			if(r_axi_wr_req == 1) begin
				if(r_m_axi_awlen == 0)
					next_w_state <= S_W_DATA_LAST;
				else
					next_w_state <= S_W_DATA;
			end
			else
				next_w_state <= S_W_IDLE;
		end
		S_W_DATA: begin
			if(m_axi_wready == 1) begin
				if(r_wr_data_cnt == 2)
					next_w_state <= S_W_DATA_LAST;
				else
					next_w_state <= S_W_DATA;
			end
			else
				next_w_state <= S_W_READY_WAIT;
		end
		S_W_READY_WAIT: begin
			if(m_axi_wready == 1) begin
				if(r_wr_data_cnt == 0)
					next_w_state <= S_W_DATA_LAST;
				else
					next_w_state <= S_W_DATA;
			end
			else
				next_w_state <= S_W_READY_WAIT;
		end
		S_W_DATA_LAST: begin
			if(m_axi_wready == 1)
				next_w_state <= S_W_IDLE;
			else
				next_w_state <= S_W_DATA_LAST;
		end
		default: begin
			next_w_state <= S_W_IDLE;
		end
	endcase
end

always @ (posedge m_axi_aclk)
begin
	case(cur_w_state)
		S_W_IDLE: begin
			r_wr_data_cnt <= r_m_axi_awlen;
			r_pcie_rx_fifo_rd_data <= pcie_rx_fifo_rd_data;
		end
		S_W_DATA: begin
			r_wr_data_cnt <= r_wr_data_cnt - 2;
			r_pcie_rx_fifo_rd_data <= pcie_rx_fifo_rd_data;
			r_pcie_rx_fifo_rd_data_d1 <= r_pcie_rx_fifo_rd_data;
		end
		S_W_READY_WAIT: begin

		end
		S_W_DATA_LAST: begin

		end
		default: begin

		end
	endcase
end

always @ (*)
begin
	if(r_m_axi_wdata_sel == 1)
		r_m_axi_wdata <= r_pcie_rx_fifo_rd_data_d1;
	else
		r_m_axi_wdata <= r_pcie_rx_fifo_rd_data;
end

always @ (*)
begin
	case(cur_w_state)
		S_W_IDLE: begin
			r_m_axi_wdata_sel <= 0;
			r_m_axi_wlast <= 0;
			r_m_axi_wvalid <= 0;
			r_axi_wr_rdy <= 1;
			r_pcie_rx_fifo_rd_en <= r_axi_wr_req;
		end
		S_W_DATA: begin
			r_m_axi_wdata_sel <= 0;
			r_m_axi_wlast <= 0;
			r_m_axi_wvalid <= 1;
			r_axi_wr_rdy <= 0;
			r_pcie_rx_fifo_rd_en <= 1;
		end
		S_W_READY_WAIT: begin
			r_m_axi_wdata_sel <= 1;
			r_m_axi_wlast <= 0;
			r_m_axi_wvalid <= 1;
			r_axi_wr_rdy <= 0;
			r_pcie_rx_fifo_rd_en <= 0;
		end
		S_W_DATA_LAST: begin
			r_m_axi_wdata_sel <= 0;
			r_m_axi_wlast <= 1;
			r_m_axi_wvalid <= 1;
			r_axi_wr_rdy <= 0;
			r_pcie_rx_fifo_rd_en <= 0;
		end
		default: begin
			r_m_axi_wdata_sel <= 0;
			r_m_axi_wlast <= 0;
			r_m_axi_wvalid <= 0;
			r_axi_wr_rdy <= 0;
			r_pcie_rx_fifo_rd_en <= 0;
		end
	endcase
end

endmodule
