

// * v1.0.0
//   - first draft
//////////////////////////////////////////////////////////////////////////////////

`define D_SC_GF_ORDER 12 // Galois field order, GF(2^12)
`define D_SC_ECC_T 14 // error correction capability t = 14

`define D_SC_P_LVL 8 // data area BCH decoder SC parallel level, 8bit I/F with NAND

`define D_SC_I_CNT 277 // received coded message length, (256B chunk + 21B parity) / 8b = 277
`define D_SC_I_CNT_BIT 9 // 2^8 = 256

`define D_SC_MSG_LENGTH 256 // message length, 256B chunk / 8b = 256
`define D_SC_MSG_LENGTH_BIT 8 // 2^8 = 256
