

`timescale 1ns / 1ps

  module dma_done # (
	parameter 	P_SLOT_TAG_WIDTH			=  10, //slot_modified
	parameter	C_PCIE_DATA_WIDTH			= 512,
	parameter	C_PCIE_ADDR_WIDTH			= 48 //modified
)
(
  	input									pcie_user_clk,
  	input									pcie_user_rst_n,

  	output									dma_done_rd_en,
  	input	[(P_SLOT_TAG_WIDTH+15)-1:0]		dma_done_rd_data, //slot_modified
  	input									dma_done_empty_n,

  	output	[P_SLOT_TAG_WIDTH-1:0]			hcmd_nlb_rd_addr, //slot_modified
  	input	[18:0]							hcmd_nlb_rd_data,

  	output									hcmd_nlb_wr1_en,
  	output	[P_SLOT_TAG_WIDTH-1:0]			hcmd_nlb_wr1_addr, //slot_modified
  	output	[18:0]							hcmd_nlb_wr1_data,
  	input									hcmd_nlb_wr1_rdy_n,

  	output									hcmd_cq_wr0_en,
  	output	[(P_SLOT_TAG_WIDTH+28)-1:0]		hcmd_cq_wr0_data0, //slot_modified
  	output	[(P_SLOT_TAG_WIDTH+28)-1:0]		hcmd_cq_wr0_data1, //slot_modified
  	input									hcmd_cq_wr0_rdy_n,

  	input									cpu_bus_clk,
  	input									cpu_bus_rst_n,

  	output	[7:0]							dma_rx_direct_done_cnt,
  	output	[7:0]							dma_tx_direct_done_cnt,
  	output	[7:0]							dma_rx_done_cnt,
  	output	[7:0]							dma_tx_done_cnt

);

localparam	LP_NLB_WR_DELAY					= 1;

localparam	S_IDLE							= 11'b00000000001;
localparam	S_DMA_INFO						= 11'b00000000010;
localparam	S_NLB_RD_WAIT					= 11'b00000000100;
localparam	S_NLB_INFO						= 11'b00000001000;
localparam	S_NLB_CALC						= 11'b00000010000;
localparam	S_NLB_WR_WAIT					= 11'b00000100000;
localparam	S_NLB_WR						= 11'b00001000000;
localparam	S_NLB_WR_DELAY					= 11'b00010000000;
localparam	S_CQ_WR_WAIT					= 11'b00100000000;
localparam	S_CQ_WR							= 11'b01000000000;
localparam	S_NLB_DONE						= 11'b10000000000;
    
      reg		[10:0]								cur_state;
      reg		[10:0]								next_state;
    
      reg											r_dma_cmd_type;
      reg											r_dma_cmd_auto_cpl;
      reg											r_dma_done_check;
      reg											r_dma_dir;
      reg		[P_SLOT_TAG_WIDTH-1:0]				r_hcmd_slot_tag; //slot_modified
      reg		[12:2]								r_dma_len;
      reg		[20:2]								r_hcmd_data_len;
    
      reg											r_dma_done_rd_en;
      reg											r_hcmd_nlb_wr1_en;
      reg											r_hcmd_cq_wr0_en;
    
      reg											r_dma_rx_direct_done_en;
      reg											r_dma_tx_direct_done_en;
      reg											r_dma_rx_done_en;
      reg											r_dma_tx_done_en;
    
      reg											r_dma_rx_direct_done_en_d1;
      reg											r_dma_tx_direct_done_en_d1;
      reg											r_dma_rx_done_en_d1;
      reg											r_dma_tx_done_en_d1;
    
      reg											r_dma_rx_direct_done_en_sync;
      reg											r_dma_tx_direct_done_en_sync;
      reg											r_dma_rx_done_en_sync;
      reg											r_dma_tx_done_en_sync;
    
      reg		[3:0]								r_nlb_wr_delay;
    
     (* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_dma_rx_direct_done;
     (* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_dma_tx_direct_done;
     (* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_dma_rx_done;
     (* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_dma_tx_done;
    
     (* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_dma_rx_direct_done_d1;
     (* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_dma_tx_direct_done_d1;
     (* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_dma_rx_done_d1;
     (* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_dma_tx_done_d1;
    
     (* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_dma_rx_direct_done_d2;
     (* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_dma_tx_direct_done_d2;
     (* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_dma_rx_done_d2;
     (* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_dma_tx_done_d2;
    
      reg		[7:0]								r_dma_rx_direct_done_cnt;
      reg		[7:0]								r_dma_tx_direct_done_cnt;
      reg		[7:0]								r_dma_rx_done_cnt;
      reg		[7:0]								r_dma_tx_done_cnt;
reg 										r_2nd_dma_need;

assign dma_done_rd_en = r_dma_done_rd_en;

assign hcmd_nlb_rd_addr = r_hcmd_slot_tag;//slot_modified

assign hcmd_nlb_wr1_en = r_hcmd_nlb_wr1_en;
assign hcmd_nlb_wr1_addr = r_hcmd_slot_tag;//slot_modified
assign hcmd_nlb_wr1_data = r_hcmd_data_len;

assign hcmd_cq_wr0_en = r_hcmd_cq_wr0_en;
assign hcmd_cq_wr0_data0 = {26'b0, r_hcmd_slot_tag, 1'b0, 1'b1}; //slot_modified
assign hcmd_cq_wr0_data1 = {(P_SLOT_TAG_WIDTH+28){1'b0}}; //slot_modified

assign dma_rx_direct_done_cnt = r_dma_rx_direct_done_cnt;
assign dma_tx_direct_done_cnt = r_dma_tx_direct_done_cnt;
assign dma_rx_done_cnt = r_dma_rx_done_cnt;
assign dma_tx_done_cnt = r_dma_tx_done_cnt;

always @ (posedge cpu_bus_clk or negedge cpu_bus_rst_n)
begin
	if(cpu_bus_rst_n == 0) begin
		r_dma_rx_direct_done_cnt <= 0;
		r_dma_tx_direct_done_cnt <= 0;
		r_dma_rx_done_cnt <= 0;
		r_dma_tx_done_cnt <= 0;
	end
	else begin
		if(r_dma_rx_direct_done_d1 == 1 && r_dma_rx_direct_done_d2 == 0)
			r_dma_rx_direct_done_cnt <= r_dma_rx_direct_done_cnt + 1;
		
		if(r_dma_tx_direct_done_d1 == 1 && r_dma_tx_direct_done_d2 == 0)
			r_dma_tx_direct_done_cnt <= r_dma_tx_direct_done_cnt + 1;

		if(r_dma_rx_done_d1 == 1 && r_dma_rx_done_d2 == 0)
			r_dma_rx_done_cnt <= r_dma_rx_done_cnt + 1;

		if(r_dma_tx_done_d1 == 1 && r_dma_tx_done_d2 == 0)
			r_dma_tx_done_cnt <= r_dma_tx_done_cnt + 1;
	end
end

always @ (posedge cpu_bus_clk)
begin
	r_dma_rx_direct_done <= r_dma_rx_direct_done_en_sync;
	r_dma_tx_direct_done <= r_dma_tx_direct_done_en_sync;
	r_dma_rx_done <= r_dma_rx_done_en_sync;
	r_dma_tx_done <= r_dma_tx_done_en_sync;

	r_dma_rx_direct_done_d1 <= r_dma_rx_direct_done;
	r_dma_tx_direct_done_d1 <= r_dma_tx_direct_done;
	r_dma_rx_done_d1 <= r_dma_rx_done;
	r_dma_tx_done_d1 <= r_dma_tx_done;

	r_dma_rx_direct_done_d2 <= r_dma_rx_direct_done_d1;
	r_dma_tx_direct_done_d2 <= r_dma_tx_direct_done_d1;
	r_dma_rx_done_d2 <= r_dma_rx_done_d1;
	r_dma_tx_done_d2 <= r_dma_tx_done_d1;
end

always @ (posedge pcie_user_clk)
begin
	r_dma_rx_direct_done_en_d1 <= r_dma_rx_direct_done_en;
	r_dma_tx_direct_done_en_d1 <= r_dma_tx_direct_done_en;
	r_dma_rx_done_en_d1 <= r_dma_rx_done_en;
	r_dma_tx_done_en_d1 <= r_dma_tx_done_en;

	r_dma_rx_direct_done_en_sync <= r_dma_rx_direct_done_en | r_dma_rx_direct_done_en_d1;
	r_dma_tx_direct_done_en_sync <= r_dma_tx_direct_done_en | r_dma_tx_direct_done_en_d1;
	r_dma_rx_done_en_sync <= r_dma_rx_done_en | r_dma_rx_done_en_d1;
	r_dma_tx_done_en_sync <= r_dma_tx_done_en | r_dma_tx_done_en_d1;
end

always @ (posedge pcie_user_clk or negedge pcie_user_rst_n)
begin
	if(pcie_user_rst_n == 0)
		cur_state <= S_IDLE;
	else
		cur_state <= next_state;
end

always @ (*)
begin
	case(cur_state)
		S_IDLE: begin
			if(dma_done_empty_n == 1'b1)
				next_state <= S_DMA_INFO;
			else
				next_state <= S_IDLE;
		end
		S_DMA_INFO: begin
			next_state <= S_NLB_RD_WAIT;
		end
		S_NLB_RD_WAIT: begin
			if(r_dma_cmd_type == 1)
				next_state <= S_NLB_DONE;
			else
				next_state <= S_NLB_INFO;
		end
		S_NLB_INFO: begin
			next_state <= S_NLB_CALC;
		end
		S_NLB_CALC: begin
            if(r_hcmd_data_len == r_dma_len) begin
                 if(r_dma_cmd_auto_cpl == 1'b1)
                     next_state <= S_CQ_WR_WAIT;
                 else
                     next_state <= S_NLB_DONE;
             end
             else
                    next_state <= S_NLB_WR_WAIT;
		end
		S_NLB_WR_WAIT: begin
			if(hcmd_nlb_wr1_rdy_n == 1)
				next_state <= S_NLB_WR_WAIT;
			else
				next_state <= S_NLB_WR;
		end
		S_NLB_WR: begin
			next_state <= S_NLB_WR_DELAY;
		end
		S_NLB_WR_DELAY: begin
			if(r_nlb_wr_delay == 0)
				next_state <= S_NLB_DONE;
			else
				next_state <= S_NLB_WR_DELAY;
		end
		S_CQ_WR_WAIT: begin
			if(hcmd_cq_wr0_rdy_n == 1)
				next_state <= S_CQ_WR_WAIT;
			else
				next_state <= S_CQ_WR;
		end
		S_CQ_WR: begin
			next_state <= S_NLB_DONE;
		end
		S_NLB_DONE: begin
			next_state <= S_IDLE;
		end
		default: begin
			next_state <= S_IDLE;
		end
	endcase
end

always @ (posedge pcie_user_clk)
begin
	case(cur_state)
		S_IDLE: begin

		end
		S_DMA_INFO: begin
		    r_dma_cmd_auto_cpl <= (r_2nd_dma_need == 1'b1 && r_dma_cmd_auto_cpl == 1'b1) ? 1'b1 : dma_done_rd_data[P_SLOT_TAG_WIDTH+14];//slot_modified
			r_dma_cmd_type <= dma_done_rd_data[P_SLOT_TAG_WIDTH+13];//slot_modified
			r_dma_done_check <= dma_done_rd_data[P_SLOT_TAG_WIDTH+12];//slot_modified
			r_dma_dir <= dma_done_rd_data[P_SLOT_TAG_WIDTH+11];//slot_modified
			r_hcmd_slot_tag <= dma_done_rd_data[(P_SLOT_TAG_WIDTH+11)-1:11]; //slot_modified
			r_dma_len <= dma_done_rd_data[10:0];
		end
		S_NLB_RD_WAIT: begin
        if(r_dma_len[11:2] != 10'b0) begin
            if(r_2nd_dma_need == 1'b1)
                r_2nd_dma_need <= 1'b0;
            else
                r_2nd_dma_need <= 1'b1;
        end
        else
            r_2nd_dma_need <= 1'b0;
		end
		S_NLB_INFO: begin
			r_hcmd_data_len <= hcmd_nlb_rd_data;
		end
		S_NLB_CALC: begin
			r_hcmd_data_len <= r_hcmd_data_len - r_dma_len;
		end
		S_NLB_WR_WAIT: begin

		end
		S_NLB_WR: begin
			r_nlb_wr_delay <= LP_NLB_WR_DELAY;
		end
		S_NLB_WR_DELAY: begin
			r_nlb_wr_delay <= r_nlb_wr_delay - 1;
		end
		S_CQ_WR_WAIT: begin

		end
		S_CQ_WR: begin

		end
		S_NLB_DONE: begin

		end
		default: begin

		end
	endcase
end

always @ (*)
begin
	case(cur_state)
		S_IDLE: begin
			r_dma_done_rd_en <= 0;
			r_hcmd_nlb_wr1_en <= 0;
			r_hcmd_cq_wr0_en <= 0;
			r_dma_rx_direct_done_en <= 0;
			r_dma_tx_direct_done_en <= 0;
			r_dma_rx_done_en <= 0;
			r_dma_tx_done_en <= 0;
		end
		S_DMA_INFO: begin
			r_dma_done_rd_en <= 1;
			r_hcmd_nlb_wr1_en <= 0;
			r_hcmd_cq_wr0_en <= 0;
			r_dma_rx_direct_done_en <= 0;
			r_dma_tx_direct_done_en <= 0;
			r_dma_rx_done_en <= 0;
			r_dma_tx_done_en <= 0;
		end
		S_NLB_RD_WAIT: begin
			r_dma_done_rd_en <= 0;
			r_hcmd_nlb_wr1_en <= 0;
			r_hcmd_cq_wr0_en <= 0;
			r_dma_rx_direct_done_en <= 0;
			r_dma_tx_direct_done_en <= 0;
			r_dma_rx_done_en <= 0;
			r_dma_tx_done_en <= 0;
		end
		S_NLB_INFO: begin
			r_dma_done_rd_en <= 0;
			r_hcmd_nlb_wr1_en <= 0;
			r_hcmd_cq_wr0_en <= 0;
			r_dma_rx_direct_done_en <= 0;
			r_dma_tx_direct_done_en <= 0;
			r_dma_rx_done_en <= 0;
			r_dma_tx_done_en <= 0;
		end
		S_NLB_CALC: begin
			r_dma_done_rd_en <= 0;
			r_hcmd_nlb_wr1_en <= 0;
			r_hcmd_cq_wr0_en <= 0;
			r_dma_rx_direct_done_en <= 0;
			r_dma_tx_direct_done_en <= 0;
			r_dma_rx_done_en <= 0;
			r_dma_tx_done_en <= 0;
		end
		S_NLB_WR_WAIT: begin
			r_dma_done_rd_en <= 0;
			r_hcmd_nlb_wr1_en <= 0;
			r_hcmd_cq_wr0_en <= 0;
			r_dma_rx_direct_done_en <= 0;
			r_dma_tx_direct_done_en <= 0;
			r_dma_rx_done_en <= 0;
			r_dma_tx_done_en <= 0;
		end
		S_NLB_WR: begin
			r_dma_done_rd_en <= 0;
			r_hcmd_nlb_wr1_en <= 1;
			r_hcmd_cq_wr0_en <= 0;
			r_dma_rx_direct_done_en <= 0;
			r_dma_tx_direct_done_en <= 0;
			r_dma_rx_done_en <= 0;
			r_dma_tx_done_en <= 0;
		end
		S_NLB_WR_DELAY: begin
			r_dma_done_rd_en <= 0;
			r_hcmd_nlb_wr1_en <= 0;
			r_hcmd_cq_wr0_en <= 0;
			r_dma_rx_direct_done_en <= 0;
			r_dma_tx_direct_done_en <= 0;
			r_dma_rx_done_en <= 0;
			r_dma_tx_done_en <= 0;
		end
		S_CQ_WR_WAIT: begin
			r_dma_done_rd_en <= 0;
			r_hcmd_nlb_wr1_en <= 0;
			r_hcmd_cq_wr0_en <= 0;
			r_dma_rx_direct_done_en <= 0;
			r_dma_tx_direct_done_en <= 0;
			r_dma_rx_done_en <= 0;
			r_dma_tx_done_en <= 0;
		end
		S_CQ_WR: begin
			r_dma_done_rd_en <= 0;
			r_hcmd_nlb_wr1_en <= 0;
			r_hcmd_cq_wr0_en <= 1;
			r_dma_rx_direct_done_en <= 0;
			r_dma_tx_direct_done_en <= 0;
			r_dma_rx_done_en <= 0;
			r_dma_tx_done_en <= 0;
		end
		S_NLB_DONE: begin
			r_dma_done_rd_en <= 0;
			r_hcmd_nlb_wr1_en <= 0;
			r_hcmd_cq_wr0_en <= 0;
			r_dma_rx_direct_done_en <= r_dma_cmd_type & r_dma_done_check & ~r_dma_dir;
			r_dma_tx_direct_done_en <= r_dma_cmd_type & r_dma_done_check & r_dma_dir;
			r_dma_rx_done_en <= ~r_dma_cmd_type & r_dma_done_check & ~r_dma_dir;
			r_dma_tx_done_en <= ~r_dma_cmd_type & r_dma_done_check & r_dma_dir;
		end
		default: begin
			r_dma_done_rd_en <= 0;
			r_hcmd_nlb_wr1_en <= 0;
			r_hcmd_cq_wr0_en <= 0;
			r_dma_rx_direct_done_en <= 0;
			r_dma_tx_direct_done_en <= 0;
			r_dma_rx_done_en <= 0;
			r_dma_tx_done_en <= 0;
		end
	endcase
end

endmodule
