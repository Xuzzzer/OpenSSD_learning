

`timescale 1ns / 1ps

module dma_cmd_fifo # (
	parameter	P_FIFO_DATA_WIDTH			= 56, //modified
	parameter	P_FIFO_DEPTH_WIDTH			= 9
)
(
	input									wr_clk,
	input									wr_rst_n,

	input									dma_cmd_wr_en,
	input	[P_FIFO_DATA_WIDTH-1:0]			dma_cmd_wr_data0,
	input	[P_FIFO_DATA_WIDTH-1:0]			dma_cmd_wr_data1,
	output									dma_cmd_wr_rdy_n,

	input									rd_clk,
	input									rd_rst_n,

	input									rd_en,
	output	[P_FIFO_DATA_WIDTH-1:0]			rd_data,
	output									empty_n
);

localparam P_FIFO_ALLOC_WIDTH				= 1;			//128 bits

localparam	S_IDLE							= 3'b001;
localparam	S_WRITE_0						= 3'b010;
localparam	S_WRITE_1						= 3'b100;

reg		[2:0]								cur_state;
reg		[2:0]								next_state;

localparam	S_SYNC_STAGE0					= 3'b001;
localparam	S_SYNC_STAGE1					= 3'b010;
localparam	S_SYNC_STAGE2					= 3'b100;

reg		[2:0]								cur_wr_state;
reg		[2:0]								next_wr_state;

reg		[2:0]								cur_rd_state;
reg		[2:0]								next_rd_state;

reg		[P_FIFO_DEPTH_WIDTH:0]				r_rear_addr;
(* KEEP = "TRUE", EQUIVALENT_REGISTER_REMOVAL = "NO" *)	reg											r_rear_sync;
(* KEEP = "TRUE", EQUIVALENT_REGISTER_REMOVAL = "NO" *)	reg											r_rear_sync_en;
reg		[P_FIFO_DEPTH_WIDTH
		:P_FIFO_ALLOC_WIDTH]				r_rear_sync_data;

(* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_front_sync_en_d1;
(* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_front_sync_en_d2;
(* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg		[P_FIFO_DEPTH_WIDTH
														:P_FIFO_ALLOC_WIDTH]				r_front_sync_addr;

reg		[P_FIFO_DEPTH_WIDTH:0]				r_front_addr;
reg		[P_FIFO_DEPTH_WIDTH:0]				r_front_addr_p1;
(* KEEP = "TRUE", EQUIVALENT_REGISTER_REMOVAL = "NO" *)	reg											r_front_sync;
(* KEEP = "TRUE", EQUIVALENT_REGISTER_REMOVAL = "NO" *)	reg											r_front_sync_en;
reg		[P_FIFO_DEPTH_WIDTH
		:P_FIFO_ALLOC_WIDTH]				r_front_sync_data;

(* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_rear_sync_en_d1;
(* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg											r_rear_sync_en_d2;
(* KEEP = "TRUE", SHIFT_EXTRACT = "NO" *)	reg		[P_FIFO_DEPTH_WIDTH
														:P_FIFO_ALLOC_WIDTH]				r_rear_sync_addr;

wire	[P_FIFO_DEPTH_WIDTH-1:0]			w_front_addr;

reg											r_wr_en;
reg											r_wr_data_sel;
reg		[P_FIFO_DATA_WIDTH-1:0]				r_wr_data;
wire										w_full_n;

reg		[P_FIFO_DATA_WIDTH-1:0]				r_dma_cmd_wr_data0;
reg		[P_FIFO_DATA_WIDTH-1:0]				r_dma_cmd_wr_data1;
reg											r_dma_cmd_wr_rdy_n;

assign dma_cmd_wr_rdy_n = r_dma_cmd_wr_rdy_n | ~w_full_n;

always @ (posedge wr_clk or negedge wr_rst_n)
begin
	if(wr_rst_n == 0)
		cur_state <= S_IDLE;
	else
		cur_state <= next_state;
end

always @ (*)
begin
	case(cur_state)
		S_IDLE: begin
			if(dma_cmd_wr_en == 1)
				next_state <= S_WRITE_0;
			else
				next_state <= S_IDLE;
		end
		S_WRITE_0: begin
			next_state <= S_WRITE_1;
		end
		S_WRITE_1: begin
			next_state <= S_IDLE;
		end
		default: begin
			next_state <= S_IDLE;
		end
	endcase
end

always @ (posedge wr_clk)
begin
	case(cur_state)
		S_IDLE: begin
			r_dma_cmd_wr_data0 <= dma_cmd_wr_data0;
			r_dma_cmd_wr_data1 <= dma_cmd_wr_data1;
		end
		S_WRITE_0: begin

		end
		S_WRITE_1: begin

		end
		default: begin

		end
	endcase
end

always @ (*)
begin
	case(cur_state)
		S_IDLE: begin
			r_wr_en <= 0;
			r_wr_data_sel <= 0;
			r_dma_cmd_wr_rdy_n <= 0;
		end
		S_WRITE_0: begin
			r_wr_en <= 1;
			r_wr_data_sel <= 0;
			r_dma_cmd_wr_rdy_n <= 1;
		end
		S_WRITE_1: begin
			r_wr_en <= 1;
			r_wr_data_sel <= 1;
			r_dma_cmd_wr_rdy_n <= 1;
		end
		default: begin
			r_wr_en <= 0;
			r_wr_data_sel <= 0;
			r_dma_cmd_wr_rdy_n <= 0;
		end
	endcase
end

always @ (*)
begin
	if(r_wr_data_sel == 0)
		r_wr_data <= r_dma_cmd_wr_data0;
	else
		r_wr_data <= r_dma_cmd_wr_data1;
end

assign w_full_n = ~((r_rear_addr[P_FIFO_DEPTH_WIDTH] ^ r_front_sync_addr[P_FIFO_DEPTH_WIDTH])
					& (r_rear_addr[P_FIFO_DEPTH_WIDTH-1:P_FIFO_ALLOC_WIDTH] 
					== r_front_sync_addr[P_FIFO_DEPTH_WIDTH-1:P_FIFO_ALLOC_WIDTH]));

always @(posedge wr_clk or negedge wr_rst_n)
begin
	if (wr_rst_n == 0) begin
		r_rear_addr <= 0;
	end
	else begin
		if (r_wr_en == 1)
			r_rear_addr  <= r_rear_addr + 1;
	end
end

assign empty_n = ~(r_front_addr[P_FIFO_DEPTH_WIDTH:P_FIFO_ALLOC_WIDTH] 
					== r_rear_sync_addr);

always @(posedge rd_clk or negedge rd_rst_n)
begin
	if (rd_rst_n == 0) begin
		r_front_addr <= 0;
		r_front_addr_p1 <= 1;
	end
	else begin
		if (rd_en == 1) begin
			r_front_addr <= r_front_addr_p1;
			r_front_addr_p1 <= r_front_addr_p1 + 1;
		end
	end
end

assign w_front_addr = (rd_en == 1) ? r_front_addr_p1[P_FIFO_DEPTH_WIDTH-1:0] 
								: r_front_addr[P_FIFO_DEPTH_WIDTH-1:0];

/////////////////////////////////////////////////////////////////////////////////////////////


always @ (posedge wr_clk or negedge wr_rst_n)
begin
	if(wr_rst_n == 0)
		cur_wr_state <= S_SYNC_STAGE0;
	else
		cur_wr_state <= next_wr_state;
end

always @(posedge wr_clk or negedge wr_rst_n)
begin
	if(wr_rst_n == 0)
		r_rear_sync_en <= 0;
	else
		r_rear_sync_en <= r_rear_sync;
end

always @(posedge wr_clk)
begin
	r_front_sync_en_d1 <= r_front_sync_en;
	r_front_sync_en_d2 <= r_front_sync_en_d1;
end

always @ (*)
begin
	case(cur_wr_state)
		S_SYNC_STAGE0: begin
			if(r_front_sync_en_d2 == 1)
				next_wr_state <= S_SYNC_STAGE1;
			else
				next_wr_state <= S_SYNC_STAGE0;
		end
		S_SYNC_STAGE1: begin
			next_wr_state <= S_SYNC_STAGE2;
		end
		S_SYNC_STAGE2: begin
			if(r_front_sync_en_d2 == 0)
				next_wr_state <= S_SYNC_STAGE0;
			else
				next_wr_state <= S_SYNC_STAGE2;
		end
		default: begin
			next_wr_state <= S_SYNC_STAGE0;
		end
	endcase
end

always @ (posedge wr_clk or negedge wr_rst_n)
begin
	if(wr_rst_n == 0) begin
		r_rear_sync_data <= 0;
		r_front_sync_addr <= 0;
	end
	else begin
		case(cur_wr_state)
			S_SYNC_STAGE0: begin

			end
			S_SYNC_STAGE1: begin
				r_rear_sync_data <= r_rear_addr[P_FIFO_DEPTH_WIDTH:P_FIFO_ALLOC_WIDTH];
				r_front_sync_addr <= r_front_sync_data;
			end
			S_SYNC_STAGE2: begin

			end
			default: begin

			end
		endcase
	end
end

always @ (*)
begin
	case(cur_wr_state)
		S_SYNC_STAGE0: begin
			r_rear_sync <= 0;
		end
		S_SYNC_STAGE1: begin
			r_rear_sync <= 0;
		end
		S_SYNC_STAGE2: begin
			r_rear_sync <= 1;
		end
		default: begin
			r_rear_sync <= 0;
		end
	endcase
end


always @ (posedge rd_clk or negedge rd_rst_n)
begin
	if(rd_rst_n == 0)
		cur_rd_state <= S_SYNC_STAGE0;
	else
		cur_rd_state <= next_rd_state;
end

always @(posedge rd_clk or negedge rd_rst_n)
begin
	if(rd_rst_n == 0)
		r_front_sync_en <= 0;
	else
		r_front_sync_en <= r_front_sync;
end

always @(posedge rd_clk)
begin
	r_rear_sync_en_d1 <= r_rear_sync_en;
	r_rear_sync_en_d2 <= r_rear_sync_en_d1;
end

always @ (*)
begin
	case(cur_rd_state)
		S_SYNC_STAGE0: begin
			if(r_rear_sync_en_d2 == 1)
				next_rd_state <= S_SYNC_STAGE1;
			else
				next_rd_state <= S_SYNC_STAGE0;
		end
		S_SYNC_STAGE1: begin
			next_rd_state <= S_SYNC_STAGE2;
		end
		S_SYNC_STAGE2: begin
			if(r_rear_sync_en_d2 == 0)
				next_rd_state <= S_SYNC_STAGE0;
			else
				next_rd_state <= S_SYNC_STAGE2;
		end
		default: begin
			next_rd_state <= S_SYNC_STAGE0;
		end
	endcase
end

always @ (posedge rd_clk or negedge rd_rst_n)
begin
	if(rd_rst_n == 0) begin
		r_front_sync_data <= 0;
		r_rear_sync_addr <= 0;
	end
	else begin
		case(cur_rd_state)
			S_SYNC_STAGE0: begin

			end
			S_SYNC_STAGE1: begin
				r_front_sync_data <= r_front_addr[P_FIFO_DEPTH_WIDTH:P_FIFO_ALLOC_WIDTH];
				r_rear_sync_addr <= r_rear_sync_data;
			end
			S_SYNC_STAGE2: begin

			end
			default: begin

			end
		endcase
	end
end

always @ (*)
begin
	case(cur_rd_state)
		S_SYNC_STAGE0: begin
			r_front_sync <= 1;
		end
		S_SYNC_STAGE1: begin
			r_front_sync <= 1;
		end
		S_SYNC_STAGE2: begin
			r_front_sync <= 0;
		end
		default: begin
			r_front_sync <= 0;
		end
	endcase
end


/////////////////////////////////////////////////////////////////////////////////////////////


localparam LP_DEVICE = "7SERIES";
localparam LP_BRAM_SIZE = "36Kb";
localparam LP_DOB_REG = 0;
localparam LP_READ_WIDTH = P_FIFO_DATA_WIDTH;
localparam LP_WRITE_WIDTH = P_FIFO_DATA_WIDTH;
localparam LP_WRITE_MODE = "WRITE_FIRST";
localparam LP_WE_WIDTH = 8;
localparam LP_ADDR_TOTAL_WITDH = 9;
localparam LP_ADDR_ZERO_PAD_WITDH = LP_ADDR_TOTAL_WITDH - P_FIFO_DEPTH_WIDTH;


generate
	wire	[LP_ADDR_TOTAL_WITDH-1:0]			rdaddr;
	wire	[LP_ADDR_TOTAL_WITDH-1:0]			wraddr;
	wire	[LP_ADDR_ZERO_PAD_WITDH-1:0]		zero_padding = 0;

	if(LP_ADDR_ZERO_PAD_WITDH == 0) begin : CALC_ADDR
		assign rdaddr = w_front_addr[P_FIFO_DEPTH_WIDTH-1:0];
		assign wraddr = r_rear_addr[P_FIFO_DEPTH_WIDTH-1:0];
	end
	else begin
		wire	[LP_ADDR_ZERO_PAD_WITDH-1:0]	zero_padding = 0;
		assign rdaddr = {zero_padding, w_front_addr[P_FIFO_DEPTH_WIDTH-1:0]};
		assign wraddr = {zero_padding, r_rear_addr[P_FIFO_DEPTH_WIDTH-1:0]};
	end
endgenerate


BRAM_SDP_MACRO #(
	.DEVICE									(LP_DEVICE),
	.BRAM_SIZE								(LP_BRAM_SIZE),
	.DO_REG									(LP_DOB_REG),
	.READ_WIDTH								(LP_READ_WIDTH),
	.WRITE_WIDTH							(LP_WRITE_WIDTH),
	.WRITE_MODE								(LP_WRITE_MODE)
)
ramb36sdp_0(
	.DO										(rd_data),
	.DI										(r_wr_data),
	.RDADDR									(rdaddr),
	.RDCLK									(rd_clk),
	.RDEN									(1'b1),
	.REGCE									(1'b1),
	.RST									(1'b0),

	.WRADDR									(wraddr),
	.WRCLK									(wr_clk),
	.WREN									(r_wr_en)
);


endmodule

