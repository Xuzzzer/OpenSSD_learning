


`define D_KES_GF_ORDER 12 // Galois field order, GF(2^15)

`define D_KES_ECC_T 14 // error correction capability t = 32
`define D_KES_ECC_T_BIT 4 // must be bigger than D_KES_ECC_T, 2^6 = 64

`define D_KES_L_CNT 14 // key equation solver loop count, D_KES_ECC_T = 32
`define D_KES_L_CNT_BIT 4 // must be bigger than D_KES_L_CNT, 2^6 = 64

//parameter ECC_PARAM_T = 32; // t = 32
//parameter KES_LOOP_COUNT = 32; // t = 32
//parameter KES_LOOP_COUNT_BIT = 6; // must be bigger than t, 2^6 = 64
